magic
tech sky130A
magscale 1 2
timestamp 1738624466
<< nwell >>
rect -38 261 2062 582
<< pwell >>
rect 12 21 2016 203
rect 29 -17 63 21
<< scnmos >>
rect 94 47 124 177
rect 178 47 208 177
rect 262 47 292 177
rect 346 47 376 177
rect 430 47 460 177
rect 514 47 544 177
rect 598 47 628 177
rect 682 47 712 177
rect 872 47 902 177
rect 956 47 986 177
rect 1040 47 1070 177
rect 1124 47 1154 177
rect 1208 47 1238 177
rect 1292 47 1322 177
rect 1376 47 1406 177
rect 1460 47 1490 177
rect 1652 47 1682 177
rect 1736 47 1766 177
rect 1820 47 1850 177
rect 1904 47 1934 177
<< scpmoshvt >>
rect 94 297 124 497
rect 178 297 208 497
rect 262 297 292 497
rect 346 297 376 497
rect 430 297 460 497
rect 514 297 544 497
rect 598 297 628 497
rect 682 297 712 497
rect 872 297 902 497
rect 956 297 986 497
rect 1040 297 1070 497
rect 1124 297 1154 497
rect 1208 297 1238 497
rect 1292 297 1322 497
rect 1376 297 1406 497
rect 1460 297 1490 497
rect 1652 297 1682 497
rect 1736 297 1766 497
rect 1820 297 1850 497
rect 1904 297 1934 497
<< ndiff >>
rect 38 95 94 177
rect 38 61 50 95
rect 84 61 94 95
rect 38 47 94 61
rect 124 163 178 177
rect 124 129 134 163
rect 168 129 178 163
rect 124 47 178 129
rect 208 95 262 177
rect 208 61 218 95
rect 252 61 262 95
rect 208 47 262 61
rect 292 163 346 177
rect 292 129 302 163
rect 336 129 346 163
rect 292 47 346 129
rect 376 163 430 177
rect 376 129 386 163
rect 420 129 430 163
rect 376 95 430 129
rect 376 61 386 95
rect 420 61 430 95
rect 376 47 430 61
rect 460 95 514 177
rect 460 61 470 95
rect 504 61 514 95
rect 460 47 514 61
rect 544 163 598 177
rect 544 129 554 163
rect 588 129 598 163
rect 544 95 598 129
rect 544 61 554 95
rect 588 61 598 95
rect 544 47 598 61
rect 628 95 682 177
rect 628 61 638 95
rect 672 61 682 95
rect 628 47 682 61
rect 712 163 764 177
rect 712 129 722 163
rect 756 129 764 163
rect 712 95 764 129
rect 712 61 722 95
rect 756 61 764 95
rect 712 47 764 61
rect 820 163 872 177
rect 820 129 828 163
rect 862 129 872 163
rect 820 95 872 129
rect 820 61 828 95
rect 862 61 872 95
rect 820 47 872 61
rect 902 163 956 177
rect 902 129 912 163
rect 946 129 956 163
rect 902 95 956 129
rect 902 61 912 95
rect 946 61 956 95
rect 902 47 956 61
rect 986 95 1040 177
rect 986 61 996 95
rect 1030 61 1040 95
rect 986 47 1040 61
rect 1070 163 1124 177
rect 1070 129 1080 163
rect 1114 129 1124 163
rect 1070 95 1124 129
rect 1070 61 1080 95
rect 1114 61 1124 95
rect 1070 47 1124 61
rect 1154 95 1208 177
rect 1154 61 1164 95
rect 1198 61 1208 95
rect 1154 47 1208 61
rect 1238 163 1292 177
rect 1238 129 1248 163
rect 1282 129 1292 163
rect 1238 95 1292 129
rect 1238 61 1248 95
rect 1282 61 1292 95
rect 1238 47 1292 61
rect 1322 95 1376 177
rect 1322 61 1332 95
rect 1366 61 1376 95
rect 1322 47 1376 61
rect 1406 163 1460 177
rect 1406 129 1416 163
rect 1450 129 1460 163
rect 1406 95 1460 129
rect 1406 61 1416 95
rect 1450 61 1460 95
rect 1406 47 1460 61
rect 1490 95 1542 177
rect 1490 61 1500 95
rect 1534 61 1542 95
rect 1490 47 1542 61
rect 1600 163 1652 177
rect 1600 129 1608 163
rect 1642 129 1652 163
rect 1600 95 1652 129
rect 1600 61 1608 95
rect 1642 61 1652 95
rect 1600 47 1652 61
rect 1682 163 1736 177
rect 1682 129 1692 163
rect 1726 129 1736 163
rect 1682 47 1736 129
rect 1766 95 1820 177
rect 1766 61 1776 95
rect 1810 61 1820 95
rect 1766 47 1820 61
rect 1850 163 1904 177
rect 1850 129 1860 163
rect 1894 129 1904 163
rect 1850 47 1904 129
rect 1934 95 1990 177
rect 1934 61 1944 95
rect 1978 61 1990 95
rect 1934 47 1990 61
<< pdiff >>
rect 38 477 94 497
rect 38 443 50 477
rect 84 443 94 477
rect 38 409 94 443
rect 38 375 50 409
rect 84 375 94 409
rect 38 341 94 375
rect 38 307 50 341
rect 84 307 94 341
rect 38 297 94 307
rect 124 485 178 497
rect 124 451 134 485
rect 168 451 178 485
rect 124 417 178 451
rect 124 383 134 417
rect 168 383 178 417
rect 124 297 178 383
rect 208 477 262 497
rect 208 443 218 477
rect 252 443 262 477
rect 208 409 262 443
rect 208 375 218 409
rect 252 375 262 409
rect 208 341 262 375
rect 208 307 218 341
rect 252 307 262 341
rect 208 297 262 307
rect 292 485 346 497
rect 292 451 302 485
rect 336 451 346 485
rect 292 297 346 451
rect 376 477 430 497
rect 376 443 386 477
rect 420 443 430 477
rect 376 409 430 443
rect 376 375 386 409
rect 420 375 430 409
rect 376 297 430 375
rect 460 485 514 497
rect 460 451 470 485
rect 504 451 514 485
rect 460 297 514 451
rect 544 477 598 497
rect 544 443 554 477
rect 588 443 598 477
rect 544 409 598 443
rect 544 375 554 409
rect 588 375 598 409
rect 544 297 598 375
rect 628 485 682 497
rect 628 451 638 485
rect 672 451 682 485
rect 628 297 682 451
rect 712 477 764 497
rect 712 443 722 477
rect 756 443 764 477
rect 712 409 764 443
rect 712 375 722 409
rect 756 375 764 409
rect 712 297 764 375
rect 820 477 872 497
rect 820 443 828 477
rect 862 443 872 477
rect 820 409 872 443
rect 820 375 828 409
rect 862 375 872 409
rect 820 297 872 375
rect 902 485 956 497
rect 902 451 912 485
rect 946 451 956 485
rect 902 297 956 451
rect 986 477 1040 497
rect 986 443 996 477
rect 1030 443 1040 477
rect 986 409 1040 443
rect 986 375 996 409
rect 1030 375 1040 409
rect 986 297 1040 375
rect 1070 485 1124 497
rect 1070 451 1080 485
rect 1114 451 1124 485
rect 1070 297 1124 451
rect 1154 477 1208 497
rect 1154 443 1164 477
rect 1198 443 1208 477
rect 1154 409 1208 443
rect 1154 375 1164 409
rect 1198 375 1208 409
rect 1154 297 1208 375
rect 1238 409 1292 497
rect 1238 375 1248 409
rect 1282 375 1292 409
rect 1238 297 1292 375
rect 1322 477 1376 497
rect 1322 443 1332 477
rect 1366 443 1376 477
rect 1322 297 1376 443
rect 1406 409 1460 497
rect 1406 375 1416 409
rect 1450 375 1460 409
rect 1406 297 1460 375
rect 1490 477 1542 497
rect 1490 443 1500 477
rect 1534 443 1542 477
rect 1490 297 1542 443
rect 1596 477 1652 497
rect 1596 443 1608 477
rect 1642 443 1652 477
rect 1596 409 1652 443
rect 1596 375 1608 409
rect 1642 375 1652 409
rect 1596 341 1652 375
rect 1596 307 1608 341
rect 1642 307 1652 341
rect 1596 297 1652 307
rect 1682 485 1736 497
rect 1682 451 1692 485
rect 1726 451 1736 485
rect 1682 417 1736 451
rect 1682 383 1692 417
rect 1726 383 1736 417
rect 1682 297 1736 383
rect 1766 477 1820 497
rect 1766 443 1776 477
rect 1810 443 1820 477
rect 1766 409 1820 443
rect 1766 375 1776 409
rect 1810 375 1820 409
rect 1766 341 1820 375
rect 1766 307 1776 341
rect 1810 307 1820 341
rect 1766 297 1820 307
rect 1850 485 1904 497
rect 1850 451 1860 485
rect 1894 451 1904 485
rect 1850 417 1904 451
rect 1850 383 1860 417
rect 1894 383 1904 417
rect 1850 297 1904 383
rect 1934 477 1990 497
rect 1934 443 1944 477
rect 1978 443 1990 477
rect 1934 409 1990 443
rect 1934 375 1944 409
rect 1978 375 1990 409
rect 1934 341 1990 375
rect 1934 307 1944 341
rect 1978 307 1990 341
rect 1934 297 1990 307
<< ndiffc >>
rect 50 61 84 95
rect 134 129 168 163
rect 218 61 252 95
rect 302 129 336 163
rect 386 129 420 163
rect 386 61 420 95
rect 470 61 504 95
rect 554 129 588 163
rect 554 61 588 95
rect 638 61 672 95
rect 722 129 756 163
rect 722 61 756 95
rect 828 129 862 163
rect 828 61 862 95
rect 912 129 946 163
rect 912 61 946 95
rect 996 61 1030 95
rect 1080 129 1114 163
rect 1080 61 1114 95
rect 1164 61 1198 95
rect 1248 129 1282 163
rect 1248 61 1282 95
rect 1332 61 1366 95
rect 1416 129 1450 163
rect 1416 61 1450 95
rect 1500 61 1534 95
rect 1608 129 1642 163
rect 1608 61 1642 95
rect 1692 129 1726 163
rect 1776 61 1810 95
rect 1860 129 1894 163
rect 1944 61 1978 95
<< pdiffc >>
rect 50 443 84 477
rect 50 375 84 409
rect 50 307 84 341
rect 134 451 168 485
rect 134 383 168 417
rect 218 443 252 477
rect 218 375 252 409
rect 218 307 252 341
rect 302 451 336 485
rect 386 443 420 477
rect 386 375 420 409
rect 470 451 504 485
rect 554 443 588 477
rect 554 375 588 409
rect 638 451 672 485
rect 722 443 756 477
rect 722 375 756 409
rect 828 443 862 477
rect 828 375 862 409
rect 912 451 946 485
rect 996 443 1030 477
rect 996 375 1030 409
rect 1080 451 1114 485
rect 1164 443 1198 477
rect 1164 375 1198 409
rect 1248 375 1282 409
rect 1332 443 1366 477
rect 1416 375 1450 409
rect 1500 443 1534 477
rect 1608 443 1642 477
rect 1608 375 1642 409
rect 1608 307 1642 341
rect 1692 451 1726 485
rect 1692 383 1726 417
rect 1776 443 1810 477
rect 1776 375 1810 409
rect 1776 307 1810 341
rect 1860 451 1894 485
rect 1860 383 1894 417
rect 1944 443 1978 477
rect 1944 375 1978 409
rect 1944 307 1978 341
<< poly >>
rect 94 497 124 523
rect 178 497 208 523
rect 262 497 292 523
rect 346 497 376 523
rect 430 497 460 523
rect 514 497 544 523
rect 598 497 628 523
rect 682 497 712 523
rect 872 497 902 523
rect 956 497 986 523
rect 1040 497 1070 523
rect 1124 497 1154 523
rect 1208 497 1238 523
rect 1292 497 1322 523
rect 1376 497 1406 523
rect 1460 497 1490 523
rect 1652 497 1682 523
rect 1736 497 1766 523
rect 1820 497 1850 523
rect 1904 497 1934 523
rect 94 265 124 297
rect 178 265 208 297
rect 262 265 292 297
rect 346 265 376 297
rect 94 249 376 265
rect 94 215 114 249
rect 148 215 182 249
rect 216 215 250 249
rect 284 215 318 249
rect 352 215 376 249
rect 94 199 376 215
rect 94 177 124 199
rect 178 177 208 199
rect 262 177 292 199
rect 346 177 376 199
rect 430 265 460 297
rect 514 265 544 297
rect 598 265 628 297
rect 682 265 712 297
rect 430 249 712 265
rect 430 215 453 249
rect 487 215 521 249
rect 555 215 589 249
rect 623 215 657 249
rect 691 215 712 249
rect 430 199 712 215
rect 430 177 460 199
rect 514 177 544 199
rect 598 177 628 199
rect 682 177 712 199
rect 872 265 902 297
rect 956 265 986 297
rect 1040 265 1070 297
rect 1124 265 1154 297
rect 872 249 1154 265
rect 872 215 892 249
rect 926 215 960 249
rect 994 215 1028 249
rect 1062 215 1154 249
rect 872 199 1154 215
rect 872 177 902 199
rect 956 177 986 199
rect 1040 177 1070 199
rect 1124 177 1154 199
rect 1208 265 1238 297
rect 1292 265 1322 297
rect 1376 265 1406 297
rect 1460 265 1490 297
rect 1208 249 1490 265
rect 1208 215 1231 249
rect 1265 215 1299 249
rect 1333 215 1367 249
rect 1401 215 1435 249
rect 1469 215 1490 249
rect 1208 199 1490 215
rect 1208 177 1238 199
rect 1292 177 1322 199
rect 1376 177 1406 199
rect 1460 177 1490 199
rect 1652 265 1682 297
rect 1736 265 1766 297
rect 1820 265 1850 297
rect 1904 265 1934 297
rect 1652 249 1934 265
rect 1652 215 1672 249
rect 1706 215 1740 249
rect 1774 215 1808 249
rect 1842 215 1876 249
rect 1910 215 1934 249
rect 1652 199 1934 215
rect 1652 177 1682 199
rect 1736 177 1766 199
rect 1820 177 1850 199
rect 1904 177 1934 199
rect 94 21 124 47
rect 178 21 208 47
rect 262 21 292 47
rect 346 21 376 47
rect 430 21 460 47
rect 514 21 544 47
rect 598 21 628 47
rect 682 21 712 47
rect 872 21 902 47
rect 956 21 986 47
rect 1040 21 1070 47
rect 1124 21 1154 47
rect 1208 21 1238 47
rect 1292 21 1322 47
rect 1376 21 1406 47
rect 1460 21 1490 47
rect 1652 21 1682 47
rect 1736 21 1766 47
rect 1820 21 1850 47
rect 1904 21 1934 47
<< polycont >>
rect 114 215 148 249
rect 182 215 216 249
rect 250 215 284 249
rect 318 215 352 249
rect 453 215 487 249
rect 521 215 555 249
rect 589 215 623 249
rect 657 215 691 249
rect 892 215 926 249
rect 960 215 994 249
rect 1028 215 1062 249
rect 1231 215 1265 249
rect 1299 215 1333 249
rect 1367 215 1401 249
rect 1435 215 1469 249
rect 1672 215 1706 249
rect 1740 215 1774 249
rect 1808 215 1842 249
rect 1876 215 1910 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 17 477 92 493
rect 17 443 50 477
rect 84 443 92 477
rect 17 409 92 443
rect 17 375 50 409
rect 84 375 92 409
rect 17 341 92 375
rect 126 485 176 527
rect 126 451 134 485
rect 168 451 176 485
rect 126 417 176 451
rect 126 383 134 417
rect 168 383 176 417
rect 126 367 176 383
rect 210 477 260 493
rect 210 443 218 477
rect 252 443 260 477
rect 210 409 260 443
rect 294 485 344 527
rect 294 451 302 485
rect 336 451 344 485
rect 294 435 344 451
rect 378 477 428 493
rect 378 443 386 477
rect 420 443 428 477
rect 210 375 218 409
rect 252 401 260 409
rect 378 409 428 443
rect 462 485 512 527
rect 462 451 470 485
rect 504 451 512 485
rect 462 435 512 451
rect 546 477 596 493
rect 546 443 554 477
rect 588 443 596 477
rect 378 401 386 409
rect 252 375 386 401
rect 420 401 428 409
rect 546 409 596 443
rect 630 485 680 527
rect 630 451 638 485
rect 672 451 680 485
rect 630 435 680 451
rect 714 477 764 493
rect 714 443 722 477
rect 756 443 764 477
rect 546 401 554 409
rect 420 375 554 401
rect 588 401 596 409
rect 714 409 764 443
rect 714 401 722 409
rect 588 375 722 401
rect 756 375 764 409
rect 17 307 50 341
rect 84 323 92 341
rect 210 357 764 375
rect 807 477 870 493
rect 807 443 828 477
rect 862 443 870 477
rect 807 409 870 443
rect 904 485 954 527
rect 904 451 912 485
rect 946 451 954 485
rect 904 435 954 451
rect 988 477 1038 493
rect 988 443 996 477
rect 1030 443 1038 477
rect 807 375 828 409
rect 862 401 870 409
rect 988 409 1038 443
rect 1072 485 1122 527
rect 1072 451 1080 485
rect 1114 451 1122 485
rect 1072 435 1122 451
rect 1156 477 1550 493
rect 1156 443 1164 477
rect 1198 443 1332 477
rect 1366 443 1500 477
rect 1534 443 1550 477
rect 1592 477 1650 493
rect 1592 443 1608 477
rect 1642 443 1650 477
rect 988 401 996 409
rect 862 375 996 401
rect 1030 401 1038 409
rect 1156 409 1198 443
rect 1592 409 1650 443
rect 1156 401 1164 409
rect 1030 375 1164 401
rect 807 357 1198 375
rect 1232 375 1248 409
rect 1282 375 1416 409
rect 1450 375 1608 409
rect 1642 375 1650 409
rect 1232 357 1650 375
rect 1684 485 1734 527
rect 1684 451 1692 485
rect 1726 451 1734 485
rect 1684 417 1734 451
rect 1684 383 1692 417
rect 1726 383 1734 417
rect 1684 367 1734 383
rect 1768 477 1818 493
rect 1768 443 1776 477
rect 1810 443 1818 477
rect 1768 409 1818 443
rect 1768 375 1776 409
rect 1810 375 1818 409
rect 210 341 260 357
rect 210 323 218 341
rect 84 307 213 323
rect 252 307 260 341
rect 1592 341 1650 357
rect 17 289 213 307
rect 247 289 260 307
rect 337 289 1146 323
rect 1180 289 1225 323
rect 1259 289 1554 323
rect 1592 307 1608 341
rect 1642 333 1650 341
rect 1768 341 1818 375
rect 1852 485 1902 527
rect 1852 451 1860 485
rect 1894 451 1902 485
rect 1852 417 1902 451
rect 1852 383 1860 417
rect 1894 383 1902 417
rect 1852 367 1902 383
rect 1936 477 2007 493
rect 1936 443 1944 477
rect 1978 443 2007 477
rect 1936 409 2007 443
rect 1936 375 1944 409
rect 1978 375 2007 409
rect 1768 333 1776 341
rect 1642 307 1776 333
rect 1810 333 1818 341
rect 1936 341 2007 375
rect 1936 333 1944 341
rect 1810 307 1944 333
rect 1978 307 2007 341
rect 1592 289 2007 307
rect 17 181 64 289
rect 337 255 371 289
rect 1112 255 1146 289
rect 1520 255 1554 289
rect 98 249 371 255
rect 98 215 114 249
rect 148 215 182 249
rect 216 215 250 249
rect 284 215 318 249
rect 352 215 371 249
rect 435 249 1078 255
rect 435 215 453 249
rect 487 215 521 249
rect 555 215 589 249
rect 623 215 657 249
rect 691 215 892 249
rect 926 215 960 249
rect 994 215 1028 249
rect 1062 215 1078 249
rect 1112 249 1486 255
rect 1112 215 1231 249
rect 1265 215 1299 249
rect 1333 215 1367 249
rect 1401 215 1435 249
rect 1469 215 1486 249
rect 1520 249 1929 255
rect 1520 215 1672 249
rect 1706 215 1740 249
rect 1774 215 1808 249
rect 1842 215 1876 249
rect 1910 215 1929 249
rect 1963 181 2007 289
rect 17 163 352 181
rect 17 129 134 163
rect 168 129 302 163
rect 336 129 352 163
rect 386 163 772 181
rect 420 145 554 163
rect 420 129 436 145
rect 386 95 436 129
rect 538 129 554 145
rect 588 145 722 163
rect 588 129 604 145
rect 34 61 50 95
rect 84 61 218 95
rect 252 61 386 95
rect 420 61 436 95
rect 34 51 436 61
rect 470 95 504 111
rect 470 17 504 61
rect 538 95 604 129
rect 706 129 722 145
rect 756 129 772 163
rect 538 61 554 95
rect 588 61 604 95
rect 538 51 604 61
rect 638 95 672 111
rect 638 17 672 61
rect 706 95 772 129
rect 706 61 722 95
rect 756 61 772 95
rect 706 51 772 61
rect 807 163 862 181
rect 807 129 828 163
rect 807 95 862 129
rect 807 61 828 95
rect 807 17 862 61
rect 896 163 1642 181
rect 896 129 912 163
rect 946 145 1080 163
rect 946 129 962 145
rect 896 95 962 129
rect 1064 129 1080 145
rect 1114 145 1248 163
rect 1114 129 1130 145
rect 896 61 912 95
rect 946 61 962 95
rect 896 51 962 61
rect 996 95 1030 111
rect 996 17 1030 61
rect 1064 95 1130 129
rect 1232 129 1248 145
rect 1282 145 1416 163
rect 1282 129 1298 145
rect 1064 61 1080 95
rect 1114 61 1130 95
rect 1064 51 1130 61
rect 1164 95 1198 111
rect 1164 17 1198 61
rect 1232 95 1298 129
rect 1400 129 1416 145
rect 1450 147 1608 163
rect 1450 145 1486 147
rect 1450 129 1466 145
rect 1232 61 1248 95
rect 1282 61 1298 95
rect 1232 51 1298 61
rect 1332 95 1366 111
rect 1332 17 1366 61
rect 1400 95 1466 129
rect 1592 129 1608 147
rect 1676 163 2007 181
rect 1676 129 1692 163
rect 1726 129 1860 163
rect 1894 129 2007 163
rect 1400 61 1416 95
rect 1450 61 1466 95
rect 1400 51 1466 61
rect 1500 95 1554 111
rect 1534 61 1554 95
rect 1592 95 1642 129
rect 1592 61 1608 95
rect 1642 61 1776 95
rect 1810 61 1944 95
rect 1978 61 1994 95
rect 1500 17 1554 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 213 307 218 323
rect 218 307 247 323
rect 213 289 247 307
rect 1225 289 1259 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 201 323 259 329
rect 201 289 213 323
rect 247 320 259 323
rect 1213 323 1271 329
rect 1213 320 1225 323
rect 247 292 1225 320
rect 247 289 259 292
rect 201 283 259 289
rect 1213 289 1225 292
rect 1259 289 1271 323
rect 1213 283 1271 289
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< labels >>
flabel locali s 1965 357 1999 391 0 FreeSans 400 0 0 0 Y
port 6 nsew
flabel locali s 213 221 247 255 0 FreeSans 400 0 0 0 B
port 7 nsew
flabel locali s 765 221 799 255 0 FreeSans 400 0 0 0 A
port 8 nsew
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 2 nsew
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 3 nsew
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
rlabel comment s 0 0 0 0 4 xnor2_4
<< properties >>
string FIXED_BBOX 0 0 2024 544
string GDS_END 378258
string GDS_FILE ./clock-divider/mag_gds/clock_divider.gds
string GDS_START 364218
string path 0.000 0.000 10.120 0.000 
<< end >>
