magic
tech sky130A
magscale 1 2
timestamp 1729294469
<< viali >>
rect 5181 23273 5215 23307
rect 7665 23273 7699 23307
rect 3341 23205 3375 23239
rect 3525 23205 3559 23239
rect 4813 23205 4847 23239
rect 11069 23205 11103 23239
rect 1777 23137 1811 23171
rect 3985 23137 4019 23171
rect 4261 23137 4295 23171
rect 4997 23137 5031 23171
rect 5365 23137 5399 23171
rect 7849 23137 7883 23171
rect 13553 23137 13587 23171
rect 16497 23137 16531 23171
rect 18337 23137 18371 23171
rect 18521 23137 18555 23171
rect 19441 23137 19475 23171
rect 22385 23137 22419 23171
rect 4721 23069 4755 23103
rect 13829 23069 13863 23103
rect 19717 23069 19751 23103
rect 22569 23069 22603 23103
rect 4077 23001 4111 23035
rect 1961 22933 1995 22967
rect 3525 22933 3559 22967
rect 3709 22933 3743 22967
rect 11345 22933 11379 22967
rect 16681 22933 16715 22967
rect 18337 22933 18371 22967
rect 7665 22729 7699 22763
rect 12081 22729 12115 22763
rect 12633 22729 12667 22763
rect 17601 22729 17635 22763
rect 17785 22729 17819 22763
rect 10517 22661 10551 22695
rect 15209 22661 15243 22695
rect 20637 22661 20671 22695
rect 3801 22593 3835 22627
rect 14013 22593 14047 22627
rect 15945 22593 15979 22627
rect 18889 22593 18923 22627
rect 20913 22593 20947 22627
rect 21373 22593 21407 22627
rect 3065 22525 3099 22559
rect 3433 22525 3467 22559
rect 3617 22525 3651 22559
rect 4077 22525 4111 22559
rect 4721 22525 4755 22559
rect 5181 22525 5215 22559
rect 7297 22525 7331 22559
rect 7665 22525 7699 22559
rect 8769 22525 8803 22559
rect 10241 22525 10275 22559
rect 11805 22525 11839 22559
rect 12541 22525 12575 22559
rect 12633 22525 12667 22559
rect 12725 22525 12759 22559
rect 12818 22525 12852 22559
rect 14105 22525 14139 22559
rect 14933 22525 14967 22559
rect 15485 22525 15519 22559
rect 17877 22525 17911 22559
rect 18061 22525 18095 22559
rect 18429 22525 18463 22559
rect 18981 22525 19015 22559
rect 19809 22525 19843 22559
rect 20361 22525 20395 22559
rect 21281 22525 21315 22559
rect 21741 22525 21775 22559
rect 8401 22457 8435 22491
rect 8585 22457 8619 22491
rect 10517 22457 10551 22491
rect 12081 22457 12115 22491
rect 15209 22457 15243 22491
rect 15669 22457 15703 22491
rect 16681 22457 16715 22491
rect 17417 22457 17451 22491
rect 20637 22457 20671 22491
rect 21925 22457 21959 22491
rect 2881 22389 2915 22423
rect 7481 22389 7515 22423
rect 10333 22389 10367 22423
rect 11897 22389 11931 22423
rect 12265 22389 12299 22423
rect 13093 22389 13127 22423
rect 13737 22389 13771 22423
rect 15025 22389 15059 22423
rect 15301 22389 15335 22423
rect 17627 22389 17661 22423
rect 18337 22389 18371 22423
rect 20453 22389 20487 22423
rect 21557 22389 21591 22423
rect 13369 22185 13403 22219
rect 15669 22185 15703 22219
rect 20111 22185 20145 22219
rect 6285 22117 6319 22151
rect 6485 22117 6519 22151
rect 7389 22117 7423 22151
rect 13521 22117 13555 22151
rect 13737 22117 13771 22151
rect 15301 22117 15335 22151
rect 15501 22117 15535 22151
rect 19901 22117 19935 22151
rect 22569 22117 22603 22151
rect 22753 22117 22787 22151
rect 4261 22049 4295 22083
rect 5089 22049 5123 22083
rect 5825 22049 5859 22083
rect 6009 22049 6043 22083
rect 6745 22049 6779 22083
rect 6837 22049 6871 22083
rect 7021 22049 7055 22083
rect 7113 22049 7147 22083
rect 7757 22049 7791 22083
rect 8033 22049 8067 22083
rect 8309 22049 8343 22083
rect 8493 22049 8527 22083
rect 8585 22049 8619 22083
rect 8677 22049 8711 22083
rect 9321 22049 9355 22083
rect 9505 22049 9539 22083
rect 10425 22049 10459 22083
rect 10518 22049 10552 22083
rect 11069 22049 11103 22083
rect 12081 22049 12115 22083
rect 12541 22049 12575 22083
rect 12909 22049 12943 22083
rect 14013 22049 14047 22083
rect 14105 22049 14139 22083
rect 15025 22049 15059 22083
rect 16129 22049 16163 22083
rect 16865 22049 16899 22083
rect 17049 22049 17083 22083
rect 17693 22049 17727 22083
rect 18153 22049 18187 22083
rect 18797 22049 18831 22083
rect 20913 22049 20947 22083
rect 21097 22049 21131 22083
rect 21649 22049 21683 22083
rect 21925 22049 21959 22083
rect 22477 22049 22511 22083
rect 8125 21981 8159 22015
rect 10333 21981 10367 22015
rect 13277 21981 13311 22015
rect 13829 21981 13863 22015
rect 15117 21981 15151 22015
rect 20361 21981 20395 22015
rect 20821 21981 20855 22015
rect 22201 21981 22235 22015
rect 22293 21981 22327 22015
rect 5181 21913 5215 21947
rect 6653 21913 6687 21947
rect 8217 21913 8251 21947
rect 8953 21913 8987 21947
rect 14657 21913 14691 21947
rect 20637 21913 20671 21947
rect 22477 21913 22511 21947
rect 5917 21845 5951 21879
rect 6469 21845 6503 21879
rect 7297 21845 7331 21879
rect 10609 21845 10643 21879
rect 13553 21845 13587 21879
rect 13921 21845 13955 21879
rect 15485 21845 15519 21879
rect 16313 21845 16347 21879
rect 17785 21845 17819 21879
rect 18337 21845 18371 21879
rect 19441 21845 19475 21879
rect 20085 21845 20119 21879
rect 20269 21845 20303 21879
rect 20913 21845 20947 21879
rect 21373 21845 21407 21879
rect 22017 21845 22051 21879
rect 22109 21845 22143 21879
rect 8217 21641 8251 21675
rect 11897 21641 11931 21675
rect 16405 21641 16439 21675
rect 17417 21641 17451 21675
rect 21189 21641 21223 21675
rect 22017 21641 22051 21675
rect 7205 21573 7239 21607
rect 9689 21573 9723 21607
rect 9873 21573 9907 21607
rect 18429 21573 18463 21607
rect 20729 21573 20763 21607
rect 20913 21573 20947 21607
rect 5181 21505 5215 21539
rect 6561 21505 6595 21539
rect 7389 21505 7423 21539
rect 7849 21505 7883 21539
rect 9321 21505 9355 21539
rect 10241 21505 10275 21539
rect 11713 21505 11747 21539
rect 12265 21505 12299 21539
rect 12725 21505 12759 21539
rect 15301 21505 15335 21539
rect 16865 21505 16899 21539
rect 21097 21505 21131 21539
rect 4629 21437 4663 21471
rect 5273 21437 5307 21471
rect 7021 21437 7055 21471
rect 7481 21437 7515 21471
rect 7941 21437 7975 21471
rect 8585 21437 8619 21471
rect 8861 21437 8895 21471
rect 8953 21437 8987 21471
rect 9137 21437 9171 21471
rect 10149 21437 10183 21471
rect 10609 21437 10643 21471
rect 10885 21437 10919 21471
rect 12173 21437 12207 21471
rect 12449 21437 12483 21471
rect 13093 21437 13127 21471
rect 13185 21437 13219 21471
rect 14565 21437 14599 21471
rect 14933 21437 14967 21471
rect 15393 21437 15427 21471
rect 16773 21437 16807 21471
rect 18153 21437 18187 21471
rect 19533 21437 19567 21471
rect 19687 21437 19721 21471
rect 21373 21437 21407 21471
rect 21465 21437 21499 21471
rect 21557 21437 21591 21471
rect 21833 21437 21867 21471
rect 3893 21369 3927 21403
rect 8220 21369 8254 21403
rect 8769 21369 8803 21403
rect 9413 21369 9447 21403
rect 12081 21369 12115 21403
rect 13553 21369 13587 21403
rect 14749 21369 14783 21403
rect 16037 21369 16071 21403
rect 16221 21369 16255 21403
rect 17233 21369 17267 21403
rect 17693 21369 17727 21403
rect 17877 21369 17911 21403
rect 18429 21369 18463 21403
rect 20453 21369 20487 21403
rect 21005 21369 21039 21403
rect 5917 21301 5951 21335
rect 6009 21301 6043 21335
rect 6377 21301 6411 21335
rect 6469 21301 6503 21335
rect 6929 21301 6963 21335
rect 8033 21301 8067 21335
rect 8401 21301 8435 21335
rect 10517 21301 10551 21335
rect 10701 21301 10735 21335
rect 11069 21301 11103 21335
rect 12633 21301 12667 21335
rect 13369 21301 13403 21335
rect 15117 21301 15151 21335
rect 15761 21301 15795 21335
rect 17141 21301 17175 21335
rect 17433 21301 17467 21335
rect 17601 21301 17635 21335
rect 18061 21301 18095 21335
rect 18245 21301 18279 21335
rect 19901 21301 19935 21335
rect 21649 21301 21683 21335
rect 7757 21097 7791 21131
rect 9965 21097 9999 21131
rect 16865 21097 16899 21131
rect 8309 21029 8343 21063
rect 9045 21029 9079 21063
rect 15485 21029 15519 21063
rect 17049 21029 17083 21063
rect 4445 20961 4479 20995
rect 4997 20961 5031 20995
rect 7205 20961 7239 20995
rect 7297 20961 7331 20995
rect 7481 20961 7515 20995
rect 7573 20961 7607 20995
rect 8217 20961 8251 20995
rect 8493 20961 8527 20995
rect 8953 20961 8987 20995
rect 9137 20961 9171 20995
rect 9229 20961 9263 20995
rect 9413 20961 9447 20995
rect 9873 20961 9907 20995
rect 10057 20961 10091 20995
rect 12265 20961 12299 20995
rect 12725 20961 12759 20995
rect 13093 20961 13127 20995
rect 13277 20961 13311 20995
rect 14749 20961 14783 20995
rect 14933 20961 14967 20995
rect 15393 20961 15427 20995
rect 15577 20961 15611 20995
rect 15761 20961 15795 20995
rect 15945 20961 15979 20995
rect 16405 20961 16439 20995
rect 16589 20961 16623 20995
rect 16773 20961 16807 20995
rect 17417 20961 17451 20995
rect 19563 20961 19597 20995
rect 19717 20961 19751 20995
rect 21649 20961 21683 20995
rect 21741 20961 21775 20995
rect 22385 20961 22419 20995
rect 12633 20893 12667 20927
rect 14105 20893 14139 20927
rect 14841 20893 14875 20927
rect 15853 20893 15887 20927
rect 17509 20893 17543 20927
rect 21465 20893 21499 20927
rect 21557 20893 21591 20927
rect 8677 20825 8711 20859
rect 17049 20825 17083 20859
rect 22109 20825 22143 20859
rect 9321 20757 9355 20791
rect 12909 20757 12943 20791
rect 16221 20757 16255 20791
rect 17785 20757 17819 20791
rect 19533 20757 19567 20791
rect 21281 20757 21315 20791
rect 21925 20757 21959 20791
rect 9229 20553 9263 20587
rect 20821 20553 20855 20587
rect 21097 20553 21131 20587
rect 21557 20553 21591 20587
rect 4721 20485 4755 20519
rect 4445 20417 4479 20451
rect 4353 20349 4387 20383
rect 4813 20349 4847 20383
rect 4997 20349 5031 20383
rect 5273 20349 5307 20383
rect 5365 20349 5399 20383
rect 5549 20349 5583 20383
rect 9229 20349 9263 20383
rect 9413 20349 9447 20383
rect 19441 20349 19475 20383
rect 19625 20349 19659 20383
rect 20545 20349 20579 20383
rect 21097 20349 21131 20383
rect 21281 20349 21315 20383
rect 4905 20281 4939 20315
rect 20637 20281 20671 20315
rect 20821 20281 20855 20315
rect 21541 20281 21575 20315
rect 21741 20281 21775 20315
rect 5733 20213 5767 20247
rect 19441 20213 19475 20247
rect 20913 20213 20947 20247
rect 21373 20213 21407 20247
rect 21281 20009 21315 20043
rect 4169 19941 4203 19975
rect 4353 19941 4387 19975
rect 4813 19941 4847 19975
rect 5365 19941 5399 19975
rect 2789 19873 2823 19907
rect 2973 19873 3007 19907
rect 3525 19873 3559 19907
rect 4537 19873 4571 19907
rect 4721 19873 4755 19907
rect 4905 19873 4939 19907
rect 5181 19873 5215 19907
rect 8493 19873 8527 19907
rect 9137 19873 9171 19907
rect 9873 19873 9907 19907
rect 11161 19873 11195 19907
rect 18889 19873 18923 19907
rect 19073 19873 19107 19907
rect 19165 19873 19199 19907
rect 20545 19873 20579 19907
rect 20637 19873 20671 19907
rect 21005 19873 21039 19907
rect 21649 19873 21683 19907
rect 2881 19805 2915 19839
rect 9781 19805 9815 19839
rect 11069 19805 11103 19839
rect 21741 19805 21775 19839
rect 10241 19737 10275 19771
rect 3157 19669 3191 19703
rect 3341 19669 3375 19703
rect 5549 19669 5583 19703
rect 7665 19669 7699 19703
rect 11529 19669 11563 19703
rect 19165 19669 19199 19703
rect 20361 19669 20395 19703
rect 21925 19669 21959 19703
rect 3893 19465 3927 19499
rect 5273 19465 5307 19499
rect 5825 19465 5859 19499
rect 6193 19465 6227 19499
rect 17049 19465 17083 19499
rect 17509 19465 17543 19499
rect 2881 19397 2915 19431
rect 3525 19397 3559 19431
rect 12357 19397 12391 19431
rect 3065 19329 3099 19363
rect 3433 19329 3467 19363
rect 3985 19329 4019 19363
rect 4905 19329 4939 19363
rect 5733 19329 5767 19363
rect 6745 19329 6779 19363
rect 7297 19329 7331 19363
rect 11897 19329 11931 19363
rect 13093 19329 13127 19363
rect 13369 19329 13403 19363
rect 15945 19329 15979 19363
rect 18153 19329 18187 19363
rect 18337 19329 18371 19363
rect 19441 19329 19475 19363
rect 2605 19261 2639 19295
rect 3341 19261 3375 19295
rect 3617 19261 3651 19295
rect 3893 19261 3927 19295
rect 4997 19261 5031 19295
rect 6009 19261 6043 19295
rect 6653 19261 6687 19295
rect 7205 19261 7239 19295
rect 10241 19261 10275 19295
rect 10701 19261 10735 19295
rect 11989 19261 12023 19295
rect 13001 19261 13035 19295
rect 16037 19261 16071 19295
rect 16497 19261 16531 19295
rect 16590 19261 16624 19295
rect 16957 19261 16991 19295
rect 17141 19261 17175 19295
rect 17877 19261 17911 19295
rect 17969 19261 18003 19295
rect 18061 19261 18095 19295
rect 18705 19261 18739 19295
rect 18981 19261 19015 19295
rect 19533 19261 19567 19295
rect 19625 19261 19659 19295
rect 19717 19261 19751 19295
rect 20361 19261 20395 19295
rect 20545 19261 20579 19295
rect 20729 19261 20763 19295
rect 21005 19261 21039 19295
rect 21097 19261 21131 19295
rect 21468 19261 21502 19295
rect 22293 19261 22327 19295
rect 22385 19261 22419 19295
rect 22569 19261 22603 19295
rect 23029 19261 23063 19295
rect 6929 19193 6963 19227
rect 16865 19193 16899 19227
rect 17325 19193 17359 19227
rect 17541 19193 17575 19227
rect 20637 19193 20671 19227
rect 3801 19125 3835 19159
rect 4261 19125 4295 19159
rect 6285 19125 6319 19159
rect 7573 19125 7607 19159
rect 16405 19125 16439 19159
rect 17693 19125 17727 19159
rect 18797 19125 18831 19159
rect 19165 19125 19199 19159
rect 19257 19125 19291 19159
rect 20913 19125 20947 19159
rect 21465 19125 21499 19159
rect 21649 19125 21683 19159
rect 3249 18921 3283 18955
rect 4261 18921 4295 18955
rect 6377 18921 6411 18955
rect 16865 18921 16899 18955
rect 17693 18921 17727 18955
rect 18429 18921 18463 18955
rect 20637 18921 20671 18955
rect 2789 18853 2823 18887
rect 4445 18853 4479 18887
rect 5641 18853 5675 18887
rect 6745 18853 6779 18887
rect 8033 18853 8067 18887
rect 17877 18853 17911 18887
rect 19156 18853 19190 18887
rect 22394 18853 22428 18887
rect 3617 18785 3651 18819
rect 3709 18785 3743 18819
rect 4169 18785 4203 18819
rect 4997 18785 5031 18819
rect 6009 18785 6043 18819
rect 6469 18785 6503 18819
rect 6653 18785 6687 18819
rect 6837 18785 6871 18819
rect 7481 18785 7515 18819
rect 7849 18785 7883 18819
rect 8861 18785 8895 18819
rect 9597 18785 9631 18819
rect 10425 18785 10459 18819
rect 10609 18785 10643 18819
rect 11437 18785 11471 18819
rect 11989 18785 12023 18819
rect 12173 18785 12207 18819
rect 12725 18785 12759 18819
rect 13001 18785 13035 18819
rect 13155 18785 13189 18819
rect 14657 18785 14691 18819
rect 16497 18785 16531 18819
rect 17233 18785 17267 18819
rect 17417 18785 17451 18819
rect 17601 18785 17635 18819
rect 18061 18785 18095 18819
rect 18245 18785 18279 18819
rect 18337 18785 18371 18819
rect 18521 18785 18555 18819
rect 20821 18785 20855 18819
rect 21005 18785 21039 18819
rect 22937 18785 22971 18819
rect 5089 18717 5123 18751
rect 5917 18717 5951 18751
rect 7573 18717 7607 18751
rect 11253 18717 11287 18751
rect 11621 18717 11655 18751
rect 12449 18717 12483 18751
rect 14565 18717 14599 18751
rect 16405 18717 16439 18751
rect 18889 18717 18923 18751
rect 21097 18717 21131 18751
rect 22661 18717 22695 18751
rect 3157 18649 3191 18683
rect 4445 18649 4479 18683
rect 7113 18649 7147 18683
rect 13369 18649 13403 18683
rect 17877 18649 17911 18683
rect 3617 18581 3651 18615
rect 3985 18581 4019 18615
rect 7021 18581 7055 18615
rect 8217 18581 8251 18615
rect 8309 18581 8343 18615
rect 10425 18581 10459 18615
rect 12357 18581 12391 18615
rect 12541 18581 12575 18615
rect 12909 18581 12943 18615
rect 15025 18581 15059 18615
rect 17417 18581 17451 18615
rect 18245 18581 18279 18615
rect 20269 18581 20303 18615
rect 21281 18581 21315 18615
rect 22845 18581 22879 18615
rect 5457 18377 5491 18411
rect 12633 18377 12667 18411
rect 19717 18377 19751 18411
rect 21005 18377 21039 18411
rect 23029 18377 23063 18411
rect 11897 18309 11931 18343
rect 12909 18309 12943 18343
rect 13001 18309 13035 18343
rect 13829 18309 13863 18343
rect 16497 18309 16531 18343
rect 3433 18241 3467 18275
rect 3893 18241 3927 18275
rect 9413 18241 9447 18275
rect 10517 18241 10551 18275
rect 11437 18241 11471 18275
rect 12817 18241 12851 18275
rect 13185 18241 13219 18275
rect 15393 18241 15427 18275
rect 17233 18241 17267 18275
rect 3525 18173 3559 18207
rect 5273 18173 5307 18207
rect 7297 18173 7331 18207
rect 7481 18173 7515 18207
rect 7573 18173 7607 18207
rect 7757 18173 7791 18207
rect 8769 18173 8803 18207
rect 9597 18173 9631 18207
rect 10057 18173 10091 18207
rect 10609 18173 10643 18207
rect 10793 18173 10827 18207
rect 11161 18173 11195 18207
rect 11529 18173 11563 18207
rect 12541 18173 12575 18207
rect 12909 18173 12943 18207
rect 13553 18173 13587 18207
rect 13921 18173 13955 18207
rect 14105 18173 14139 18207
rect 15301 18173 15335 18207
rect 15761 18173 15795 18207
rect 15945 18173 15979 18207
rect 16221 18173 16255 18207
rect 16313 18173 16347 18207
rect 17417 18173 17451 18207
rect 19901 18173 19935 18207
rect 20085 18173 20119 18207
rect 20913 18173 20947 18207
rect 21649 18173 21683 18207
rect 21905 18173 21939 18207
rect 5089 18105 5123 18139
rect 8677 18105 8711 18139
rect 10333 18105 10367 18139
rect 12817 18105 12851 18139
rect 13829 18105 13863 18139
rect 16129 18105 16163 18139
rect 16497 18105 16531 18139
rect 7389 18037 7423 18071
rect 7757 18037 7791 18071
rect 11253 18037 11287 18071
rect 13645 18037 13679 18071
rect 14013 18037 14047 18071
rect 15669 18037 15703 18071
rect 17601 18037 17635 18071
rect 4261 17833 4295 17867
rect 10425 17833 10459 17867
rect 14105 17833 14139 17867
rect 21833 17765 21867 17799
rect 3617 17697 3651 17731
rect 3801 17697 3835 17731
rect 4077 17697 4111 17731
rect 9597 17697 9631 17731
rect 10057 17697 10091 17731
rect 10241 17697 10275 17731
rect 13093 17697 13127 17731
rect 13185 17697 13219 17731
rect 13737 17697 13771 17731
rect 14473 17697 14507 17731
rect 17693 17697 17727 17731
rect 17877 17697 17911 17731
rect 21649 17697 21683 17731
rect 21925 17697 21959 17731
rect 9505 17629 9539 17663
rect 9965 17629 9999 17663
rect 13645 17629 13679 17663
rect 14197 17629 14231 17663
rect 14657 17561 14691 17595
rect 13093 17493 13127 17527
rect 13461 17493 13495 17527
rect 14289 17493 14323 17527
rect 17693 17493 17727 17527
rect 21649 17493 21683 17527
rect 3893 17289 3927 17323
rect 8861 17289 8895 17323
rect 22845 17289 22879 17323
rect 18245 17221 18279 17255
rect 19073 17221 19107 17255
rect 8493 17153 8527 17187
rect 13645 17153 13679 17187
rect 14105 17153 14139 17187
rect 15669 17153 15703 17187
rect 18429 17153 18463 17187
rect 19993 17153 20027 17187
rect 5917 17085 5951 17119
rect 6101 17085 6135 17119
rect 8585 17085 8619 17119
rect 13737 17085 13771 17119
rect 15853 17085 15887 17119
rect 17877 17085 17911 17119
rect 18061 17085 18095 17119
rect 18153 17085 18187 17119
rect 18889 17085 18923 17119
rect 18981 17085 19015 17119
rect 19165 17085 19199 17119
rect 19901 17085 19935 17119
rect 20177 17085 20211 17119
rect 20453 17085 20487 17119
rect 22753 17085 22787 17119
rect 3709 17017 3743 17051
rect 18429 17017 18463 17051
rect 20361 17017 20395 17051
rect 20698 17017 20732 17051
rect 22201 17017 22235 17051
rect 22569 17017 22603 17051
rect 3909 16949 3943 16983
rect 4077 16949 4111 16983
rect 6009 16949 6043 16983
rect 16037 16949 16071 16983
rect 17969 16949 18003 16983
rect 18705 16949 18739 16983
rect 21833 16949 21867 16983
rect 3709 16745 3743 16779
rect 4261 16745 4295 16779
rect 7665 16745 7699 16779
rect 11529 16745 11563 16779
rect 18153 16745 18187 16779
rect 18613 16745 18647 16779
rect 20085 16745 20119 16779
rect 22845 16745 22879 16779
rect 2973 16677 3007 16711
rect 7297 16677 7331 16711
rect 8217 16677 8251 16711
rect 8417 16677 8451 16711
rect 12633 16677 12667 16711
rect 12817 16677 12851 16711
rect 14013 16677 14047 16711
rect 2881 16609 2915 16643
rect 3157 16609 3191 16643
rect 3341 16609 3375 16643
rect 3433 16609 3467 16643
rect 3525 16609 3559 16643
rect 3801 16609 3835 16643
rect 3985 16609 4019 16643
rect 4353 16609 4387 16643
rect 4537 16609 4571 16643
rect 4905 16609 4939 16643
rect 5549 16609 5583 16643
rect 6285 16609 6319 16643
rect 7205 16609 7239 16643
rect 7481 16609 7515 16643
rect 10425 16609 10459 16643
rect 11391 16609 11425 16643
rect 11529 16609 11563 16643
rect 11989 16609 12023 16643
rect 12449 16609 12483 16643
rect 13737 16609 13771 16643
rect 13829 16609 13863 16643
rect 15117 16609 15151 16643
rect 15301 16609 15335 16643
rect 15577 16609 15611 16643
rect 16129 16609 16163 16643
rect 16313 16609 16347 16643
rect 16589 16609 16623 16643
rect 17141 16609 17175 16643
rect 17325 16609 17359 16643
rect 17509 16609 17543 16643
rect 17785 16609 17819 16643
rect 18061 16609 18095 16643
rect 18245 16609 18279 16643
rect 18429 16609 18463 16643
rect 18972 16609 19006 16643
rect 21465 16609 21499 16643
rect 21732 16609 21766 16643
rect 6469 16541 6503 16575
rect 7021 16541 7055 16575
rect 10517 16541 10551 16575
rect 10977 16541 11011 16575
rect 12081 16541 12115 16575
rect 12357 16541 12391 16575
rect 15485 16541 15519 16575
rect 16773 16541 16807 16575
rect 18705 16541 18739 16575
rect 10793 16473 10827 16507
rect 14013 16473 14047 16507
rect 15117 16473 15151 16507
rect 8401 16405 8435 16439
rect 8585 16405 8619 16439
rect 15853 16405 15887 16439
rect 9689 16201 9723 16235
rect 9873 16201 9907 16235
rect 13553 16201 13587 16235
rect 15853 16201 15887 16235
rect 16221 16201 16255 16235
rect 16865 16201 16899 16235
rect 17049 16201 17083 16235
rect 18245 16201 18279 16235
rect 19257 16201 19291 16235
rect 21925 16201 21959 16235
rect 22017 16201 22051 16235
rect 3525 16133 3559 16167
rect 4997 16133 5031 16167
rect 8217 16133 8251 16167
rect 11437 16133 11471 16167
rect 14473 16133 14507 16167
rect 15393 16133 15427 16167
rect 16405 16133 16439 16167
rect 18107 16133 18141 16167
rect 19533 16133 19567 16167
rect 3893 16065 3927 16099
rect 4537 16065 4571 16099
rect 5917 16065 5951 16099
rect 6193 16065 6227 16099
rect 7113 16065 7147 16099
rect 7757 16065 7791 16099
rect 9229 16065 9263 16099
rect 14565 16065 14599 16099
rect 15669 16065 15703 16099
rect 21741 16065 21775 16099
rect 21833 16065 21867 16099
rect 2697 15997 2731 16031
rect 3801 15997 3835 16031
rect 4077 15997 4111 16031
rect 4629 15997 4663 16031
rect 5825 15997 5859 16031
rect 6285 15997 6319 16031
rect 6469 15997 6503 16031
rect 7205 15997 7239 16031
rect 7849 15997 7883 16031
rect 8585 15997 8619 16031
rect 8861 15997 8895 16031
rect 9045 15997 9079 16031
rect 9321 15997 9355 16031
rect 9781 15997 9815 16031
rect 9965 15997 9999 16031
rect 11161 15997 11195 16031
rect 13185 15997 13219 16031
rect 13369 15997 13403 16031
rect 13737 15997 13771 16031
rect 13921 15997 13955 16031
rect 15945 15997 15979 16031
rect 16497 15997 16531 16031
rect 16773 15997 16807 16031
rect 17049 15997 17083 16031
rect 17141 15997 17175 16031
rect 17969 15997 18003 16031
rect 18429 15997 18463 16031
rect 18705 15997 18739 16031
rect 18889 15997 18923 16031
rect 19073 15997 19107 16031
rect 19349 15997 19383 16031
rect 21465 15997 21499 16031
rect 21557 15997 21591 16031
rect 22109 15997 22143 16031
rect 2881 15929 2915 15963
rect 3249 15929 3283 15963
rect 11253 15929 11287 15963
rect 11437 15929 11471 15963
rect 14197 15929 14231 15963
rect 14657 15929 14691 15963
rect 16037 15929 16071 15963
rect 16253 15929 16287 15963
rect 16589 15929 16623 15963
rect 18981 15929 19015 15963
rect 3065 15861 3099 15895
rect 4169 15861 4203 15895
rect 6377 15861 6411 15895
rect 7573 15861 7607 15895
rect 8401 15861 8435 15895
rect 13277 15861 13311 15895
rect 14289 15861 14323 15895
rect 17417 15861 17451 15895
rect 18429 15861 18463 15895
rect 21741 15861 21775 15895
rect 3341 15657 3375 15691
rect 8033 15657 8067 15691
rect 11621 15657 11655 15691
rect 13553 15657 13587 15691
rect 22569 15657 22603 15691
rect 3683 15589 3717 15623
rect 3801 15589 3835 15623
rect 4261 15589 4295 15623
rect 4353 15589 4387 15623
rect 8585 15589 8619 15623
rect 3433 15521 3467 15555
rect 3893 15521 3927 15555
rect 3985 15521 4019 15555
rect 4629 15521 4663 15555
rect 4813 15521 4847 15555
rect 7757 15521 7791 15555
rect 7941 15521 7975 15555
rect 8309 15521 8343 15555
rect 8401 15521 8435 15555
rect 11345 15521 11379 15555
rect 11805 15521 11839 15555
rect 11897 15521 11931 15555
rect 13277 15521 13311 15555
rect 13737 15521 13771 15555
rect 13921 15521 13955 15555
rect 14013 15521 14047 15555
rect 14105 15521 14139 15555
rect 14289 15521 14323 15555
rect 15025 15521 15059 15555
rect 15209 15521 15243 15555
rect 15301 15521 15335 15555
rect 15577 15521 15611 15555
rect 18512 15521 18546 15555
rect 21741 15521 21775 15555
rect 22201 15521 22235 15555
rect 2973 15453 3007 15487
rect 3525 15453 3559 15487
rect 10977 15453 11011 15487
rect 11253 15453 11287 15487
rect 13369 15453 13403 15487
rect 14197 15453 14231 15487
rect 15117 15453 15151 15487
rect 15853 15453 15887 15487
rect 18245 15453 18279 15487
rect 21833 15453 21867 15487
rect 22293 15453 22327 15487
rect 3157 15385 3191 15419
rect 8217 15385 8251 15419
rect 12909 15385 12943 15419
rect 15485 15385 15519 15419
rect 22109 15385 22143 15419
rect 4169 15317 4203 15351
rect 8585 15317 8619 15351
rect 15669 15317 15703 15351
rect 15761 15317 15795 15351
rect 19625 15317 19659 15351
rect 22293 15317 22327 15351
rect 6009 15113 6043 15147
rect 13921 15113 13955 15147
rect 18797 15113 18831 15147
rect 4537 15045 4571 15079
rect 16589 15045 16623 15079
rect 4261 14977 4295 15011
rect 4721 14977 4755 15011
rect 5825 14977 5859 15011
rect 10885 14977 10919 15011
rect 16221 14977 16255 15011
rect 20269 14977 20303 15011
rect 21281 14977 21315 15011
rect 21557 14977 21591 15011
rect 4169 14909 4203 14943
rect 4813 14909 4847 14943
rect 5733 14909 5767 14943
rect 10977 14909 11011 14943
rect 12633 14909 12667 14943
rect 13093 14909 13127 14943
rect 13737 14909 13771 14943
rect 16037 14909 16071 14943
rect 16129 14909 16163 14943
rect 16313 14909 16347 14943
rect 16589 14909 16623 14943
rect 16773 14909 16807 14943
rect 16865 14909 16899 14943
rect 18705 14909 18739 14943
rect 18889 14909 18923 14943
rect 21189 14909 21223 14943
rect 22017 14909 22051 14943
rect 13553 14841 13587 14875
rect 19901 14841 19935 14875
rect 20085 14841 20119 14875
rect 21833 14841 21867 14875
rect 22201 14841 22235 14875
rect 5181 14773 5215 14807
rect 5365 14773 5399 14807
rect 11345 14773 11379 14807
rect 12265 14773 12299 14807
rect 16497 14773 16531 14807
rect 3065 14569 3099 14603
rect 4537 14569 4571 14603
rect 15761 14501 15795 14535
rect 19717 14501 19751 14535
rect 2697 14433 2731 14467
rect 2881 14433 2915 14467
rect 4353 14433 4387 14467
rect 4537 14433 4571 14467
rect 5181 14433 5215 14467
rect 6009 14433 6043 14467
rect 8033 14433 8067 14467
rect 9229 14433 9263 14467
rect 9322 14433 9356 14467
rect 15577 14433 15611 14467
rect 15669 14433 15703 14467
rect 15945 14433 15979 14467
rect 16129 14433 16163 14467
rect 16405 14433 16439 14467
rect 16497 14433 16531 14467
rect 18981 14433 19015 14467
rect 19165 14433 19199 14467
rect 19441 14433 19475 14467
rect 19533 14433 19567 14467
rect 19809 14433 19843 14467
rect 19993 14433 20027 14467
rect 20177 14433 20211 14467
rect 20361 14433 20395 14467
rect 20453 14433 20487 14467
rect 20545 14433 20579 14467
rect 20729 14433 20763 14467
rect 5273 14365 5307 14399
rect 5917 14365 5951 14399
rect 8125 14365 8159 14399
rect 19717 14365 19751 14399
rect 5549 14297 5583 14331
rect 9597 14297 9631 14331
rect 16221 14297 16255 14331
rect 19349 14297 19383 14331
rect 6285 14229 6319 14263
rect 8309 14229 8343 14263
rect 15393 14229 15427 14263
rect 16681 14229 16715 14263
rect 19165 14229 19199 14263
rect 19901 14229 19935 14263
rect 20177 14229 20211 14263
rect 20637 14229 20671 14263
rect 7021 14025 7055 14059
rect 8033 14025 8067 14059
rect 10701 14025 10735 14059
rect 11989 14025 12023 14059
rect 14105 14025 14139 14059
rect 16681 14025 16715 14059
rect 18153 14025 18187 14059
rect 20177 14025 20211 14059
rect 20637 14025 20671 14059
rect 20913 14025 20947 14059
rect 22661 14025 22695 14059
rect 3065 13957 3099 13991
rect 5549 13957 5583 13991
rect 6469 13957 6503 13991
rect 20729 13957 20763 13991
rect 21925 13957 21959 13991
rect 22201 13957 22235 13991
rect 5273 13889 5307 13923
rect 6009 13889 6043 13923
rect 6653 13889 6687 13923
rect 8953 13889 8987 13923
rect 9781 13889 9815 13923
rect 18705 13889 18739 13923
rect 18981 13889 19015 13923
rect 19625 13889 19659 13923
rect 19901 13889 19935 13923
rect 20269 13889 20303 13923
rect 21465 13889 21499 13923
rect 22017 13889 22051 13923
rect 22569 13889 22603 13923
rect 2789 13821 2823 13855
rect 2881 13821 2915 13855
rect 3249 13821 3283 13855
rect 3433 13821 3467 13855
rect 3617 13821 3651 13855
rect 6101 13821 6135 13855
rect 6745 13821 6779 13855
rect 7205 13821 7239 13855
rect 7298 13821 7332 13855
rect 8063 13821 8097 13855
rect 8217 13821 8251 13855
rect 9045 13821 9079 13855
rect 9689 13821 9723 13855
rect 10609 13821 10643 13855
rect 10793 13821 10827 13855
rect 11253 13821 11287 13855
rect 11345 13821 11379 13855
rect 11529 13821 11563 13855
rect 13553 13821 13587 13855
rect 13645 13821 13679 13855
rect 13829 13821 13863 13855
rect 13921 13821 13955 13855
rect 15301 13821 15335 13855
rect 15557 13821 15591 13855
rect 16773 13821 16807 13855
rect 17029 13821 17063 13855
rect 19073 13821 19107 13855
rect 19533 13821 19567 13855
rect 20453 13821 20487 13855
rect 21557 13821 21591 13855
rect 22109 13821 22143 13855
rect 22385 13821 22419 13855
rect 22477 13821 22511 13855
rect 22753 13821 22787 13855
rect 22845 13821 22879 13855
rect 20867 13787 20901 13821
rect 3065 13753 3099 13787
rect 3525 13753 3559 13787
rect 7573 13753 7607 13787
rect 11805 13753 11839 13787
rect 12005 13753 12039 13787
rect 20177 13753 20211 13787
rect 21097 13753 21131 13787
rect 3801 13685 3835 13719
rect 5733 13685 5767 13719
rect 8677 13685 8711 13719
rect 10057 13685 10091 13719
rect 11713 13685 11747 13719
rect 12173 13685 12207 13719
rect 10057 13481 10091 13515
rect 10701 13481 10735 13515
rect 12541 13481 12575 13515
rect 14473 13481 14507 13515
rect 4086 13413 4120 13447
rect 6285 13413 6319 13447
rect 9505 13413 9539 13447
rect 9721 13413 9755 13447
rect 13981 13413 14015 13447
rect 14197 13413 14231 13447
rect 17509 13413 17543 13447
rect 22687 13413 22721 13447
rect 6009 13345 6043 13379
rect 6101 13345 6135 13379
rect 9965 13345 9999 13379
rect 10241 13345 10275 13379
rect 10517 13345 10551 13379
rect 10793 13345 10827 13379
rect 12449 13345 12483 13379
rect 12725 13345 12759 13379
rect 12817 13345 12851 13379
rect 12909 13345 12943 13379
rect 13185 13345 13219 13379
rect 13277 13345 13311 13379
rect 13369 13345 13403 13379
rect 13553 13345 13587 13379
rect 14289 13345 14323 13379
rect 14565 13345 14599 13379
rect 17325 13345 17359 13379
rect 21465 13345 21499 13379
rect 21925 13345 21959 13379
rect 22201 13345 22235 13379
rect 22385 13345 22419 13379
rect 22477 13345 22511 13379
rect 22569 13345 22603 13379
rect 4353 13277 4387 13311
rect 21741 13277 21775 13311
rect 22845 13277 22879 13311
rect 6285 13209 6319 13243
rect 9873 13209 9907 13243
rect 22109 13209 22143 13243
rect 2973 13141 3007 13175
rect 9689 13141 9723 13175
rect 10425 13141 10459 13175
rect 10517 13141 10551 13175
rect 13737 13141 13771 13175
rect 13829 13141 13863 13175
rect 14013 13141 14047 13175
rect 14289 13141 14323 13175
rect 17693 13141 17727 13175
rect 21925 13141 21959 13175
rect 8769 12937 8803 12971
rect 12817 12937 12851 12971
rect 13737 12937 13771 12971
rect 17693 12937 17727 12971
rect 18245 12937 18279 12971
rect 18429 12937 18463 12971
rect 21741 12937 21775 12971
rect 9137 12869 9171 12903
rect 5181 12801 5215 12835
rect 6929 12801 6963 12835
rect 7205 12801 7239 12835
rect 8769 12801 8803 12835
rect 12081 12801 12115 12835
rect 12173 12801 12207 12835
rect 13553 12801 13587 12835
rect 15393 12801 15427 12835
rect 15485 12801 15519 12835
rect 18061 12801 18095 12835
rect 4905 12733 4939 12767
rect 6837 12733 6871 12767
rect 7297 12733 7331 12767
rect 7390 12733 7424 12767
rect 8493 12733 8527 12767
rect 8953 12733 8987 12767
rect 9229 12733 9263 12767
rect 9413 12733 9447 12767
rect 11897 12733 11931 12767
rect 11989 12733 12023 12767
rect 12357 12733 12391 12767
rect 12449 12733 12483 12767
rect 12633 12733 12667 12767
rect 12909 12733 12943 12767
rect 13002 12733 13036 12767
rect 13829 12733 13863 12767
rect 17233 12733 17267 12767
rect 17417 12733 17451 12767
rect 18245 12733 18279 12767
rect 22017 12733 22051 12767
rect 15301 12665 15335 12699
rect 17509 12665 17543 12699
rect 17969 12665 18003 12699
rect 21741 12665 21775 12699
rect 21925 12665 21959 12699
rect 4537 12597 4571 12631
rect 4997 12597 5031 12631
rect 7665 12597 7699 12631
rect 9413 12597 9447 12631
rect 11713 12597 11747 12631
rect 13277 12597 13311 12631
rect 13553 12597 13587 12631
rect 14933 12597 14967 12631
rect 17417 12597 17451 12631
rect 17709 12597 17743 12631
rect 17877 12597 17911 12631
rect 3433 12393 3467 12427
rect 5365 12393 5399 12427
rect 10349 12393 10383 12427
rect 12449 12393 12483 12427
rect 17785 12393 17819 12427
rect 18061 12393 18095 12427
rect 19073 12393 19107 12427
rect 22845 12393 22879 12427
rect 4252 12325 4286 12359
rect 8677 12325 8711 12359
rect 8861 12325 8895 12359
rect 9689 12325 9723 12359
rect 9781 12325 9815 12359
rect 10149 12325 10183 12359
rect 14832 12325 14866 12359
rect 16681 12325 16715 12359
rect 16897 12325 16931 12359
rect 17417 12325 17451 12359
rect 17969 12325 18003 12359
rect 18889 12325 18923 12359
rect 20269 12325 20303 12359
rect 20469 12325 20503 12359
rect 3985 12257 4019 12291
rect 7297 12257 7331 12291
rect 7481 12257 7515 12291
rect 8033 12257 8067 12291
rect 8217 12257 8251 12291
rect 8493 12257 8527 12291
rect 9045 12257 9079 12291
rect 9597 12257 9631 12291
rect 9965 12257 9999 12291
rect 10057 12257 10091 12291
rect 12357 12257 12391 12291
rect 12541 12257 12575 12291
rect 13277 12257 13311 12291
rect 13369 12257 13403 12291
rect 13461 12257 13495 12291
rect 17141 12257 17175 12291
rect 17233 12257 17267 12291
rect 17693 12257 17727 12291
rect 18429 12257 18463 12291
rect 18705 12257 18739 12291
rect 20729 12257 20763 12291
rect 20913 12257 20947 12291
rect 21741 12257 21775 12291
rect 21833 12257 21867 12291
rect 22293 12257 22327 12291
rect 23029 12257 23063 12291
rect 3249 12189 3283 12223
rect 3341 12189 3375 12223
rect 8125 12189 8159 12223
rect 13553 12189 13587 12223
rect 14565 12189 14599 12223
rect 18521 12189 18555 12223
rect 7481 12121 7515 12155
rect 9413 12121 9447 12155
rect 17969 12121 18003 12155
rect 22109 12121 22143 12155
rect 3801 12053 3835 12087
rect 8309 12053 8343 12087
rect 9229 12053 9263 12087
rect 10333 12053 10367 12087
rect 10517 12053 10551 12087
rect 13093 12053 13127 12087
rect 15945 12053 15979 12087
rect 16865 12053 16899 12087
rect 17049 12053 17083 12087
rect 17417 12053 17451 12087
rect 20453 12053 20487 12087
rect 20637 12053 20671 12087
rect 22017 12053 22051 12087
rect 3249 11849 3283 11883
rect 10149 11849 10183 11883
rect 16221 11849 16255 11883
rect 16405 11849 16439 11883
rect 16681 11849 16715 11883
rect 17693 11849 17727 11883
rect 19533 11849 19567 11883
rect 20085 11849 20119 11883
rect 21649 11849 21683 11883
rect 7021 11781 7055 11815
rect 20177 11781 20211 11815
rect 4629 11713 4663 11747
rect 5181 11713 5215 11747
rect 5273 11713 5307 11747
rect 10333 11713 10367 11747
rect 10701 11713 10735 11747
rect 14933 11713 14967 11747
rect 16773 11713 16807 11747
rect 21557 11713 21591 11747
rect 4362 11645 4396 11679
rect 7205 11645 7239 11679
rect 7297 11645 7331 11679
rect 7941 11645 7975 11679
rect 8125 11645 8159 11679
rect 8401 11645 8435 11679
rect 9321 11645 9355 11679
rect 9413 11645 9447 11679
rect 10057 11645 10091 11679
rect 10609 11645 10643 11679
rect 10793 11645 10827 11679
rect 10885 11645 10919 11679
rect 14666 11645 14700 11679
rect 16037 11645 16071 11679
rect 16129 11645 16163 11679
rect 16497 11645 16531 11679
rect 16589 11645 16623 11679
rect 17325 11645 17359 11679
rect 17509 11645 17543 11679
rect 19441 11645 19475 11679
rect 19625 11645 19659 11679
rect 19901 11645 19935 11679
rect 21290 11645 21324 11679
rect 23029 11645 23063 11679
rect 7021 11577 7055 11611
rect 8585 11577 8619 11611
rect 10333 11577 10367 11611
rect 19717 11577 19751 11611
rect 22762 11577 22796 11611
rect 4721 11509 4755 11543
rect 5089 11509 5123 11543
rect 8033 11509 8067 11543
rect 8769 11509 8803 11543
rect 9137 11509 9171 11543
rect 10425 11509 10459 11543
rect 13553 11509 13587 11543
rect 4629 11305 4663 11339
rect 6285 11305 6319 11339
rect 10793 11305 10827 11339
rect 11345 11305 11379 11339
rect 13553 11305 13587 11339
rect 18445 11305 18479 11339
rect 21833 11305 21867 11339
rect 3516 11237 3550 11271
rect 18245 11237 18279 11271
rect 19901 11237 19935 11271
rect 21649 11237 21683 11271
rect 22017 11237 22051 11271
rect 6193 11169 6227 11203
rect 8033 11169 8067 11203
rect 8217 11169 8251 11203
rect 10517 11169 10551 11203
rect 10609 11169 10643 11203
rect 11253 11169 11287 11203
rect 11713 11169 11747 11203
rect 11805 11169 11839 11203
rect 13737 11169 13771 11203
rect 15577 11169 15611 11203
rect 19441 11169 19475 11203
rect 20085 11169 20119 11203
rect 20821 11169 20855 11203
rect 3249 11101 3283 11135
rect 6377 11101 6411 11135
rect 13921 11101 13955 11135
rect 15669 11101 15703 11135
rect 19257 11101 19291 11135
rect 20545 11101 20579 11135
rect 20637 11101 20671 11135
rect 20729 11101 20763 11135
rect 21281 11033 21315 11067
rect 22201 11033 22235 11067
rect 5825 10965 5859 10999
rect 8125 10965 8159 10999
rect 11621 10965 11655 10999
rect 15945 10965 15979 10999
rect 18429 10965 18463 10999
rect 18613 10965 18647 10999
rect 19625 10965 19659 10999
rect 19717 10965 19751 10999
rect 21005 10965 21039 10999
rect 21649 10965 21683 10999
rect 6745 10761 6779 10795
rect 8493 10761 8527 10795
rect 10977 10761 11011 10795
rect 12449 10761 12483 10795
rect 18889 10761 18923 10795
rect 19349 10761 19383 10795
rect 21005 10761 21039 10795
rect 19257 10693 19291 10727
rect 21189 10693 21223 10727
rect 7941 10625 7975 10659
rect 8861 10625 8895 10659
rect 9045 10625 9079 10659
rect 14105 10625 14139 10659
rect 14289 10625 14323 10659
rect 5365 10557 5399 10591
rect 5632 10557 5666 10591
rect 7205 10557 7239 10591
rect 7573 10557 7607 10591
rect 7849 10557 7883 10591
rect 8401 10557 8435 10591
rect 8677 10557 8711 10591
rect 9137 10557 9171 10591
rect 9597 10557 9631 10591
rect 9864 10557 9898 10591
rect 11069 10557 11103 10591
rect 11336 10557 11370 10591
rect 18521 10557 18555 10591
rect 20729 10557 20763 10591
rect 7297 10489 7331 10523
rect 7389 10489 7423 10523
rect 18276 10489 18310 10523
rect 20462 10489 20496 10523
rect 20821 10489 20855 10523
rect 7021 10421 7055 10455
rect 8217 10421 8251 10455
rect 9505 10421 9539 10455
rect 13645 10421 13679 10455
rect 14013 10421 14047 10455
rect 17141 10421 17175 10455
rect 18705 10421 18739 10455
rect 18889 10421 18923 10455
rect 21021 10421 21055 10455
rect 4721 10217 4755 10251
rect 7941 10217 7975 10251
rect 8125 10217 8159 10251
rect 16681 10217 16715 10251
rect 17233 10217 17267 10251
rect 18153 10217 18187 10251
rect 18521 10217 18555 10251
rect 20085 10217 20119 10251
rect 22083 10217 22117 10251
rect 6828 10149 6862 10183
rect 13860 10149 13894 10183
rect 14197 10149 14231 10183
rect 15577 10149 15611 10183
rect 15777 10149 15811 10183
rect 19901 10149 19935 10183
rect 21465 10149 21499 10183
rect 22293 10149 22327 10183
rect 22569 10149 22603 10183
rect 3341 10081 3375 10115
rect 4353 10081 4387 10115
rect 4813 10081 4847 10115
rect 6561 10081 6595 10115
rect 8033 10081 8067 10115
rect 14105 10081 14139 10115
rect 14381 10081 14415 10115
rect 14565 10081 14599 10115
rect 16313 10081 16347 10115
rect 16773 10081 16807 10115
rect 17049 10081 17083 10115
rect 18061 10081 18095 10115
rect 18337 10081 18371 10115
rect 19533 10081 19567 10115
rect 22385 10081 22419 10115
rect 3433 10013 3467 10047
rect 4445 10013 4479 10047
rect 5089 10013 5123 10047
rect 14657 10013 14691 10047
rect 16221 10013 16255 10047
rect 16865 10013 16899 10047
rect 4997 9945 5031 9979
rect 21833 9945 21867 9979
rect 22753 9945 22787 9979
rect 3709 9877 3743 9911
rect 4353 9877 4387 9911
rect 4905 9877 4939 9911
rect 12725 9877 12759 9911
rect 15761 9877 15795 9911
rect 15945 9877 15979 9911
rect 16773 9877 16807 9911
rect 19901 9877 19935 9911
rect 21281 9877 21315 9911
rect 21465 9877 21499 9911
rect 21925 9877 21959 9911
rect 22109 9877 22143 9911
rect 4629 9673 4663 9707
rect 13047 9673 13081 9707
rect 14933 9673 14967 9707
rect 17417 9673 17451 9707
rect 19349 9673 19383 9707
rect 20821 9673 20855 9707
rect 21281 9673 21315 9707
rect 22753 9673 22787 9707
rect 5273 9605 5307 9639
rect 15853 9605 15887 9639
rect 18429 9605 18463 9639
rect 4721 9537 4755 9571
rect 8861 9537 8895 9571
rect 9045 9537 9079 9571
rect 10517 9537 10551 9571
rect 10701 9537 10735 9571
rect 20453 9537 20487 9571
rect 21373 9537 21407 9571
rect 4629 9469 4663 9503
rect 4905 9469 4939 9503
rect 5457 9469 5491 9503
rect 5549 9469 5583 9503
rect 5641 9469 5675 9503
rect 5825 9469 5859 9503
rect 12909 9469 12943 9503
rect 13185 9469 13219 9503
rect 13369 9469 13403 9503
rect 13553 9469 13587 9503
rect 13820 9469 13854 9503
rect 15577 9469 15611 9503
rect 15853 9469 15887 9503
rect 16405 9469 16439 9503
rect 16589 9469 16623 9503
rect 16681 9469 16715 9503
rect 16957 9469 16991 9503
rect 17049 9469 17083 9503
rect 18337 9469 18371 9503
rect 18521 9469 18555 9503
rect 18889 9469 18923 9503
rect 20637 9469 20671 9503
rect 20913 9469 20947 9503
rect 5273 9401 5307 9435
rect 13277 9401 13311 9435
rect 17417 9401 17451 9435
rect 18705 9401 18739 9435
rect 19073 9401 19107 9435
rect 19317 9401 19351 9435
rect 19533 9401 19567 9435
rect 21097 9401 21131 9435
rect 21618 9401 21652 9435
rect 5089 9333 5123 9367
rect 5825 9333 5859 9367
rect 8401 9333 8435 9367
rect 8769 9333 8803 9367
rect 10057 9333 10091 9367
rect 10425 9333 10459 9367
rect 15669 9333 15703 9367
rect 16773 9333 16807 9367
rect 17601 9333 17635 9367
rect 19165 9333 19199 9367
rect 9137 9129 9171 9163
rect 10793 9129 10827 9163
rect 14565 9129 14599 9163
rect 15945 9129 15979 9163
rect 18153 9129 18187 9163
rect 22661 9129 22695 9163
rect 3525 9061 3559 9095
rect 8024 9061 8058 9095
rect 9680 9061 9714 9095
rect 19266 9061 19300 9095
rect 3065 8993 3099 9027
rect 3249 8993 3283 9027
rect 3341 8993 3375 9027
rect 3985 8993 4019 9027
rect 4629 8993 4663 9027
rect 5089 8993 5123 9027
rect 7757 8993 7791 9027
rect 9413 8993 9447 9027
rect 11437 8993 11471 9027
rect 11713 8993 11747 9027
rect 14105 8993 14139 9027
rect 14381 8993 14415 9027
rect 15577 8993 15611 9027
rect 15761 8993 15795 9027
rect 17518 8993 17552 9027
rect 19533 8993 19567 9027
rect 21537 8993 21571 9027
rect 4077 8925 4111 8959
rect 4905 8925 4939 8959
rect 11529 8925 11563 8959
rect 14197 8925 14231 8959
rect 17785 8925 17819 8959
rect 21281 8925 21315 8959
rect 4353 8857 4387 8891
rect 16405 8857 16439 8891
rect 3157 8789 3191 8823
rect 3709 8789 3743 8823
rect 5089 8789 5123 8823
rect 5273 8789 5307 8823
rect 11437 8789 11471 8823
rect 11897 8789 11931 8823
rect 14197 8789 14231 8823
rect 3893 8585 3927 8619
rect 4813 8585 4847 8619
rect 4997 8585 5031 8619
rect 6009 8585 6043 8619
rect 7481 8585 7515 8619
rect 7757 8585 7791 8619
rect 8401 8585 8435 8619
rect 11299 8585 11333 8619
rect 15485 8585 15519 8619
rect 17141 8585 17175 8619
rect 21281 8585 21315 8619
rect 21465 8585 21499 8619
rect 6561 8517 6595 8551
rect 10609 8517 10643 8551
rect 15669 8517 15703 8551
rect 21833 8517 21867 8551
rect 7665 8449 7699 8483
rect 8585 8449 8619 8483
rect 10701 8449 10735 8483
rect 11529 8449 11563 8483
rect 13277 8449 13311 8483
rect 13645 8449 13679 8483
rect 14565 8449 14599 8483
rect 6285 8381 6319 8415
rect 6377 8381 6411 8415
rect 6561 8381 6595 8415
rect 7389 8381 7423 8415
rect 7757 8381 7791 8415
rect 7941 8381 7975 8415
rect 8677 8381 8711 8415
rect 10425 8381 10459 8415
rect 10609 8381 10643 8415
rect 10885 8381 10919 8415
rect 11161 8381 11195 8415
rect 11437 8381 11471 8415
rect 11621 8381 11655 8415
rect 12357 8381 12391 8415
rect 12541 8381 12575 8415
rect 13185 8381 13219 8415
rect 13369 8381 13403 8415
rect 13737 8381 13771 8415
rect 14381 8381 14415 8415
rect 15117 8381 15151 8415
rect 15761 8381 15795 8415
rect 16017 8381 16051 8415
rect 3939 8347 3973 8381
rect 3709 8313 3743 8347
rect 4629 8313 4663 8347
rect 4829 8313 4863 8347
rect 5825 8313 5859 8347
rect 6041 8313 6075 8347
rect 8401 8313 8435 8347
rect 14197 8313 14231 8347
rect 21465 8313 21499 8347
rect 4077 8245 4111 8279
rect 6193 8245 6227 8279
rect 7665 8245 7699 8279
rect 8125 8245 8159 8279
rect 8861 8245 8895 8279
rect 11069 8245 11103 8279
rect 12541 8245 12575 8279
rect 14105 8245 14139 8279
rect 15485 8245 15519 8279
rect 3985 8041 4019 8075
rect 4077 8041 4111 8075
rect 6285 8041 6319 8075
rect 16129 8041 16163 8075
rect 16681 8041 16715 8075
rect 16849 8041 16883 8075
rect 21281 8041 21315 8075
rect 2697 7973 2731 8007
rect 3801 7973 3835 8007
rect 7849 7973 7883 8007
rect 16497 7973 16531 8007
rect 17049 7973 17083 8007
rect 22109 7973 22143 8007
rect 2237 7905 2271 7939
rect 2421 7905 2455 7939
rect 2881 7905 2915 7939
rect 3157 7905 3191 7939
rect 3341 7905 3375 7939
rect 3433 7905 3467 7939
rect 4169 7905 4203 7939
rect 5917 7905 5951 7939
rect 6101 7905 6135 7939
rect 6561 7905 6595 7939
rect 8125 7905 8159 7939
rect 8585 7905 8619 7939
rect 11345 7905 11379 7939
rect 11621 7905 11655 7939
rect 11805 7905 11839 7939
rect 13553 7905 13587 7939
rect 13737 7905 13771 7939
rect 14013 7905 14047 7939
rect 14289 7905 14323 7939
rect 16313 7905 16347 7939
rect 16589 7905 16623 7939
rect 18705 7905 18739 7939
rect 18961 7905 18995 7939
rect 21649 7905 21683 7939
rect 21925 7905 21959 7939
rect 6469 7837 6503 7871
rect 7941 7837 7975 7871
rect 8493 7837 8527 7871
rect 11253 7837 11287 7871
rect 14105 7837 14139 7871
rect 21465 7837 21499 7871
rect 21557 7837 21591 7871
rect 21741 7837 21775 7871
rect 8953 7769 8987 7803
rect 20085 7769 20119 7803
rect 2329 7701 2363 7735
rect 2513 7701 2547 7735
rect 2973 7701 3007 7735
rect 4353 7701 4387 7735
rect 6101 7701 6135 7735
rect 6929 7701 6963 7735
rect 7941 7701 7975 7735
rect 8309 7701 8343 7735
rect 11069 7701 11103 7735
rect 11621 7701 11655 7735
rect 13737 7701 13771 7735
rect 14013 7701 14047 7735
rect 14473 7701 14507 7735
rect 16865 7701 16899 7735
rect 22293 7701 22327 7735
rect 4629 7497 4663 7531
rect 7389 7497 7423 7531
rect 7941 7497 7975 7531
rect 8401 7497 8435 7531
rect 8585 7497 8619 7531
rect 13277 7497 13311 7531
rect 14013 7497 14047 7531
rect 14289 7497 14323 7531
rect 18797 7497 18831 7531
rect 18981 7497 19015 7531
rect 19257 7497 19291 7531
rect 20729 7497 20763 7531
rect 21373 7497 21407 7531
rect 3249 7361 3283 7395
rect 7021 7361 7055 7395
rect 10793 7361 10827 7395
rect 12817 7361 12851 7395
rect 13645 7361 13679 7395
rect 14473 7361 14507 7395
rect 22201 7361 22235 7395
rect 1685 7293 1719 7327
rect 4905 7293 4939 7327
rect 7113 7293 7147 7327
rect 8125 7293 8159 7327
rect 8217 7293 8251 7327
rect 10701 7293 10735 7327
rect 12909 7293 12943 7327
rect 13737 7293 13771 7327
rect 14565 7293 14599 7327
rect 16037 7293 16071 7327
rect 16221 7293 16255 7327
rect 18337 7293 18371 7327
rect 18521 7293 18555 7327
rect 19625 7293 19659 7327
rect 20085 7293 20119 7327
rect 21005 7293 21039 7327
rect 22477 7293 22511 7327
rect 1952 7225 1986 7259
rect 3494 7225 3528 7259
rect 4721 7225 4755 7259
rect 7941 7225 7975 7259
rect 8769 7225 8803 7259
rect 18429 7225 18463 7259
rect 18949 7225 18983 7259
rect 19165 7225 19199 7259
rect 19441 7225 19475 7259
rect 19901 7225 19935 7259
rect 20713 7225 20747 7259
rect 20913 7225 20947 7259
rect 3065 7157 3099 7191
rect 5089 7157 5123 7191
rect 8559 7157 8593 7191
rect 11069 7157 11103 7191
rect 16221 7157 16255 7191
rect 19717 7157 19751 7191
rect 20545 7157 20579 7191
rect 21373 7157 21407 7191
rect 21557 7157 21591 7191
rect 2145 6953 2179 6987
rect 2313 6953 2347 6987
rect 3157 6953 3191 6987
rect 3249 6953 3283 6987
rect 4261 6953 4295 6987
rect 17509 6953 17543 6987
rect 21005 6953 21039 6987
rect 2513 6885 2547 6919
rect 2973 6885 3007 6919
rect 3417 6885 3451 6919
rect 3617 6885 3651 6919
rect 15577 6885 15611 6919
rect 15761 6885 15795 6919
rect 20821 6885 20855 6919
rect 21710 6885 21744 6919
rect 2605 6817 2639 6851
rect 5374 6817 5408 6851
rect 9597 6817 9631 6851
rect 11161 6817 11195 6851
rect 11621 6817 11655 6851
rect 11897 6817 11931 6851
rect 16396 6817 16430 6851
rect 18337 6817 18371 6851
rect 18604 6817 18638 6851
rect 19901 6817 19935 6851
rect 20085 6817 20119 6851
rect 20177 6817 20211 6851
rect 20637 6817 20671 6851
rect 20729 6817 20763 6851
rect 21465 6817 21499 6851
rect 5641 6749 5675 6783
rect 9505 6749 9539 6783
rect 11069 6749 11103 6783
rect 11713 6749 11747 6783
rect 16129 6749 16163 6783
rect 9965 6681 9999 6715
rect 11529 6681 11563 6715
rect 12081 6681 12115 6715
rect 19717 6681 19751 6715
rect 20453 6681 20487 6715
rect 2329 6613 2363 6647
rect 2973 6613 3007 6647
rect 3433 6613 3467 6647
rect 11621 6613 11655 6647
rect 15945 6613 15979 6647
rect 20177 6613 20211 6647
rect 20361 6613 20395 6647
rect 22845 6613 22879 6647
rect 4629 6409 4663 6443
rect 4813 6409 4847 6443
rect 5733 6409 5767 6443
rect 6101 6409 6135 6443
rect 6469 6409 6503 6443
rect 6929 6409 6963 6443
rect 13829 6409 13863 6443
rect 14657 6409 14691 6443
rect 16221 6409 16255 6443
rect 16405 6409 16439 6443
rect 18705 6409 18739 6443
rect 18889 6409 18923 6443
rect 19349 6409 19383 6443
rect 19809 6409 19843 6443
rect 19993 6409 20027 6443
rect 21150 6409 21184 6443
rect 4261 6341 4295 6375
rect 19257 6273 19291 6307
rect 19717 6273 19751 6307
rect 20821 6273 20855 6307
rect 6009 6205 6043 6239
rect 6193 6205 6227 6239
rect 6837 6205 6871 6239
rect 7113 6205 7147 6239
rect 7297 6205 7331 6239
rect 7389 6205 7423 6239
rect 7665 6205 7699 6239
rect 14381 6205 14415 6239
rect 19533 6205 19567 6239
rect 20729 6205 20763 6239
rect 21465 6205 21499 6239
rect 5917 6137 5951 6171
rect 7481 6137 7515 6171
rect 13645 6137 13679 6171
rect 14105 6137 14139 6171
rect 14749 6137 14783 6171
rect 14933 6137 14967 6171
rect 16037 6137 16071 6171
rect 16237 6137 16271 6171
rect 18889 6137 18923 6171
rect 19977 6137 20011 6171
rect 20177 6137 20211 6171
rect 20545 6137 20579 6171
rect 21189 6137 21223 6171
rect 21710 6137 21744 6171
rect 4629 6069 4663 6103
rect 5549 6069 5583 6103
rect 5717 6069 5751 6103
rect 6285 6069 6319 6103
rect 6469 6069 6503 6103
rect 7849 6069 7883 6103
rect 13845 6069 13879 6103
rect 14013 6069 14047 6103
rect 14289 6069 14323 6103
rect 14473 6069 14507 6103
rect 15117 6069 15151 6103
rect 21373 6069 21407 6103
rect 22845 6069 22879 6103
rect 5641 5865 5675 5899
rect 7481 5865 7515 5899
rect 7573 5865 7607 5899
rect 11253 5865 11287 5899
rect 11989 5865 12023 5899
rect 14473 5865 14507 5899
rect 19993 5865 20027 5899
rect 20453 5865 20487 5899
rect 21741 5865 21775 5899
rect 22569 5865 22603 5899
rect 5273 5797 5307 5831
rect 5457 5797 5491 5831
rect 10241 5797 10275 5831
rect 10977 5797 11011 5831
rect 11345 5797 11379 5831
rect 13645 5797 13679 5831
rect 15209 5797 15243 5831
rect 22201 5797 22235 5831
rect 6368 5729 6402 5763
rect 8686 5729 8720 5763
rect 8953 5729 8987 5763
rect 9137 5729 9171 5763
rect 9321 5729 9355 5763
rect 9873 5729 9907 5763
rect 10149 5729 10183 5763
rect 10425 5729 10459 5763
rect 11161 5729 11195 5763
rect 13001 5729 13035 5763
rect 13185 5729 13219 5763
rect 14013 5729 14047 5763
rect 14289 5729 14323 5763
rect 14565 5729 14599 5763
rect 14841 5729 14875 5763
rect 18613 5729 18647 5763
rect 18880 5729 18914 5763
rect 20269 5729 20303 5763
rect 20545 5729 20579 5763
rect 21281 5729 21315 5763
rect 21465 5729 21499 5763
rect 21925 5729 21959 5763
rect 22017 5729 22051 5763
rect 22385 5729 22419 5763
rect 6101 5661 6135 5695
rect 11529 5661 11563 5695
rect 11621 5661 11655 5695
rect 10057 5593 10091 5627
rect 13461 5593 13495 5627
rect 21649 5593 21683 5627
rect 9229 5525 9263 5559
rect 10609 5525 10643 5559
rect 11989 5525 12023 5559
rect 12173 5525 12207 5559
rect 13093 5525 13127 5559
rect 13645 5525 13679 5559
rect 14105 5525 14139 5559
rect 15209 5525 15243 5559
rect 15393 5525 15427 5559
rect 20085 5525 20119 5559
rect 21465 5525 21499 5559
rect 2697 5321 2731 5355
rect 3525 5321 3559 5355
rect 6837 5321 6871 5355
rect 8033 5321 8067 5355
rect 8217 5321 8251 5355
rect 8769 5321 8803 5355
rect 10885 5321 10919 5355
rect 10977 5321 11011 5355
rect 12725 5321 12759 5355
rect 15117 5321 15151 5355
rect 18797 5321 18831 5355
rect 18981 5321 19015 5355
rect 21741 5321 21775 5355
rect 3065 5253 3099 5287
rect 7021 5253 7055 5287
rect 7573 5253 7607 5287
rect 19349 5253 19383 5287
rect 9505 5185 9539 5219
rect 16497 5185 16531 5219
rect 5457 5117 5491 5151
rect 5713 5117 5747 5151
rect 7205 5117 7239 5151
rect 7297 5117 7331 5151
rect 7665 5117 7699 5151
rect 9413 5117 9447 5151
rect 12090 5117 12124 5151
rect 12357 5117 12391 5151
rect 13185 5117 13219 5151
rect 13369 5117 13403 5151
rect 13553 5117 13587 5151
rect 13820 5117 13854 5151
rect 16230 5117 16264 5151
rect 20269 5117 20303 5151
rect 20361 5117 20395 5151
rect 20453 5117 20487 5151
rect 20637 5117 20671 5151
rect 20729 5117 20763 5151
rect 20913 5117 20947 5151
rect 21925 5117 21959 5151
rect 3341 5049 3375 5083
rect 8033 5049 8067 5083
rect 8585 5049 8619 5083
rect 8801 5049 8835 5083
rect 9045 5049 9079 5083
rect 9229 5049 9263 5083
rect 9772 5049 9806 5083
rect 12541 5049 12575 5083
rect 12757 5049 12791 5083
rect 13001 5049 13035 5083
rect 18981 5049 19015 5083
rect 2513 4981 2547 5015
rect 2697 4981 2731 5015
rect 3541 4981 3575 5015
rect 3709 4981 3743 5015
rect 7389 4981 7423 5015
rect 8953 4981 8987 5015
rect 12909 4981 12943 5015
rect 14933 4981 14967 5015
rect 19993 4981 20027 5015
rect 20821 4981 20855 5015
rect 3801 4777 3835 4811
rect 4169 4777 4203 4811
rect 6561 4777 6595 4811
rect 8033 4777 8067 4811
rect 10149 4777 10183 4811
rect 10333 4777 10367 4811
rect 14197 4777 14231 4811
rect 21097 4777 21131 4811
rect 2666 4709 2700 4743
rect 3893 4709 3927 4743
rect 4705 4709 4739 4743
rect 4905 4709 4939 4743
rect 6193 4709 6227 4743
rect 6729 4709 6763 4743
rect 6929 4709 6963 4743
rect 8125 4709 8159 4743
rect 8944 4709 8978 4743
rect 13062 4709 13096 4743
rect 19984 4709 20018 4743
rect 2421 4641 2455 4675
rect 4077 4641 4111 4675
rect 4261 4641 4295 4675
rect 6377 4641 6411 4675
rect 11529 4641 11563 4675
rect 11805 4641 11839 4675
rect 2329 4573 2363 4607
rect 8677 4573 8711 4607
rect 12817 4573 12851 4607
rect 19717 4573 19751 4607
rect 2053 4505 2087 4539
rect 4445 4505 4479 4539
rect 10701 4505 10735 4539
rect 1869 4437 1903 4471
rect 4537 4437 4571 4471
rect 4721 4437 4755 4471
rect 6745 4437 6779 4471
rect 10057 4437 10091 4471
rect 10333 4437 10367 4471
rect 3065 4233 3099 4267
rect 10241 4233 10275 4267
rect 10425 4233 10459 4267
rect 22845 4233 22879 4267
rect 1685 4097 1719 4131
rect 3249 4097 3283 4131
rect 3617 4097 3651 4131
rect 3709 4097 3743 4131
rect 5641 4097 5675 4131
rect 11345 4097 11379 4131
rect 1941 4029 1975 4063
rect 3433 4029 3467 4063
rect 3525 4029 3559 4063
rect 4077 4029 4111 4063
rect 4344 4029 4378 4063
rect 5549 4029 5583 4063
rect 5733 4029 5767 4063
rect 10977 4029 11011 4063
rect 11161 4029 11195 4063
rect 23029 4029 23063 4063
rect 10609 3961 10643 3995
rect 5457 3893 5491 3927
rect 10399 3893 10433 3927
rect 3065 3689 3099 3723
rect 4629 3689 4663 3723
rect 4721 3689 4755 3723
rect 2973 3621 3007 3655
rect 3157 3621 3191 3655
rect 3516 3621 3550 3655
rect 5089 3621 5123 3655
rect 2881 3553 2915 3587
rect 3249 3553 3283 3587
rect 4905 3553 4939 3587
rect 3433 3145 3467 3179
rect 3617 2941 3651 2975
rect 3801 2941 3835 2975
rect 3893 2941 3927 2975
<< metal1 >>
rect 552 23418 23368 23440
rect 552 23366 4322 23418
rect 4374 23366 4386 23418
rect 4438 23366 4450 23418
rect 4502 23366 4514 23418
rect 4566 23366 4578 23418
rect 4630 23366 23368 23418
rect 552 23344 23368 23366
rect 5169 23307 5227 23313
rect 5169 23304 5181 23307
rect 3436 23276 5181 23304
rect 3436 23248 3464 23276
rect 5169 23273 5181 23276
rect 5215 23273 5227 23307
rect 5169 23267 5227 23273
rect 5258 23264 5264 23316
rect 5316 23304 5322 23316
rect 7653 23307 7711 23313
rect 7653 23304 7665 23307
rect 5316 23276 7665 23304
rect 5316 23264 5322 23276
rect 7653 23273 7665 23276
rect 7699 23273 7711 23307
rect 7653 23267 7711 23273
rect 3329 23239 3387 23245
rect 3329 23205 3341 23239
rect 3375 23236 3387 23239
rect 3418 23236 3424 23248
rect 3375 23208 3424 23236
rect 3375 23205 3387 23208
rect 3329 23199 3387 23205
rect 3418 23196 3424 23208
rect 3476 23196 3482 23248
rect 3513 23239 3571 23245
rect 3513 23205 3525 23239
rect 3559 23236 3571 23239
rect 4801 23239 4859 23245
rect 4801 23236 4813 23239
rect 3559 23208 4813 23236
rect 3559 23205 3571 23208
rect 3513 23199 3571 23205
rect 1762 23128 1768 23180
rect 1820 23128 1826 23180
rect 2774 23128 2780 23180
rect 2832 23168 2838 23180
rect 3528 23168 3556 23199
rect 3988 23177 4016 23208
rect 4801 23205 4813 23208
rect 4847 23205 4859 23239
rect 4801 23199 4859 23205
rect 4890 23196 4896 23248
rect 4948 23236 4954 23248
rect 4948 23208 5396 23236
rect 4948 23196 4954 23208
rect 2832 23140 3556 23168
rect 3973 23171 4031 23177
rect 2832 23128 2838 23140
rect 3973 23137 3985 23171
rect 4019 23137 4031 23171
rect 3973 23131 4031 23137
rect 4249 23171 4307 23177
rect 4249 23137 4261 23171
rect 4295 23137 4307 23171
rect 4249 23131 4307 23137
rect 3418 23060 3424 23112
rect 3476 23100 3482 23112
rect 4264 23100 4292 23131
rect 4338 23128 4344 23180
rect 4396 23168 4402 23180
rect 4982 23168 4988 23180
rect 4396 23140 4988 23168
rect 4396 23128 4402 23140
rect 4982 23128 4988 23140
rect 5040 23168 5046 23180
rect 5258 23168 5264 23180
rect 5040 23140 5264 23168
rect 5040 23128 5046 23140
rect 5258 23128 5264 23140
rect 5316 23128 5322 23180
rect 5368 23177 5396 23208
rect 10502 23196 10508 23248
rect 10560 23236 10566 23248
rect 11057 23239 11115 23245
rect 11057 23236 11069 23239
rect 10560 23208 11069 23236
rect 10560 23196 10566 23208
rect 11057 23205 11069 23208
rect 11103 23205 11115 23239
rect 11057 23199 11115 23205
rect 5353 23171 5411 23177
rect 5353 23137 5365 23171
rect 5399 23137 5411 23171
rect 5353 23131 5411 23137
rect 7558 23128 7564 23180
rect 7616 23168 7622 23180
rect 7837 23171 7895 23177
rect 7837 23168 7849 23171
rect 7616 23140 7849 23168
rect 7616 23128 7622 23140
rect 7837 23137 7849 23140
rect 7883 23137 7895 23171
rect 7837 23131 7895 23137
rect 13538 23128 13544 23180
rect 13596 23128 13602 23180
rect 16482 23128 16488 23180
rect 16540 23128 16546 23180
rect 17954 23128 17960 23180
rect 18012 23168 18018 23180
rect 18325 23171 18383 23177
rect 18325 23168 18337 23171
rect 18012 23140 18337 23168
rect 18012 23128 18018 23140
rect 18325 23137 18337 23140
rect 18371 23137 18383 23171
rect 18325 23131 18383 23137
rect 18509 23171 18567 23177
rect 18509 23137 18521 23171
rect 18555 23168 18567 23171
rect 18782 23168 18788 23180
rect 18555 23140 18788 23168
rect 18555 23137 18567 23140
rect 18509 23131 18567 23137
rect 18782 23128 18788 23140
rect 18840 23128 18846 23180
rect 19426 23128 19432 23180
rect 19484 23128 19490 23180
rect 22278 23128 22284 23180
rect 22336 23168 22342 23180
rect 22373 23171 22431 23177
rect 22373 23168 22385 23171
rect 22336 23140 22385 23168
rect 22336 23128 22342 23140
rect 22373 23137 22385 23140
rect 22419 23137 22431 23171
rect 22373 23131 22431 23137
rect 3476 23072 4292 23100
rect 4709 23103 4767 23109
rect 3476 23060 3482 23072
rect 4709 23069 4721 23103
rect 4755 23100 4767 23103
rect 5810 23100 5816 23112
rect 4755 23072 5816 23100
rect 4755 23069 4767 23072
rect 4709 23063 4767 23069
rect 5810 23060 5816 23072
rect 5868 23060 5874 23112
rect 13817 23103 13875 23109
rect 13817 23069 13829 23103
rect 13863 23100 13875 23103
rect 13906 23100 13912 23112
rect 13863 23072 13912 23100
rect 13863 23069 13875 23072
rect 13817 23063 13875 23069
rect 13906 23060 13912 23072
rect 13964 23060 13970 23112
rect 15194 23060 15200 23112
rect 15252 23100 15258 23112
rect 15470 23100 15476 23112
rect 15252 23072 15476 23100
rect 15252 23060 15258 23072
rect 15470 23060 15476 23072
rect 15528 23100 15534 23112
rect 18414 23100 18420 23112
rect 15528 23072 18420 23100
rect 15528 23060 15534 23072
rect 18414 23060 18420 23072
rect 18472 23100 18478 23112
rect 19705 23103 19763 23109
rect 19705 23100 19717 23103
rect 18472 23072 19717 23100
rect 18472 23060 18478 23072
rect 19705 23069 19717 23072
rect 19751 23100 19763 23103
rect 21910 23100 21916 23112
rect 19751 23072 21916 23100
rect 19751 23069 19763 23072
rect 19705 23063 19763 23069
rect 21910 23060 21916 23072
rect 21968 23060 21974 23112
rect 22002 23060 22008 23112
rect 22060 23100 22066 23112
rect 22557 23103 22615 23109
rect 22557 23100 22569 23103
rect 22060 23072 22569 23100
rect 22060 23060 22066 23072
rect 22557 23069 22569 23072
rect 22603 23069 22615 23103
rect 22557 23063 22615 23069
rect 2866 22992 2872 23044
rect 2924 23032 2930 23044
rect 4065 23035 4123 23041
rect 4065 23032 4077 23035
rect 2924 23004 4077 23032
rect 2924 22992 2930 23004
rect 1949 22967 2007 22973
rect 1949 22933 1961 22967
rect 1995 22964 2007 22967
rect 3050 22964 3056 22976
rect 1995 22936 3056 22964
rect 1995 22933 2007 22936
rect 1949 22927 2007 22933
rect 3050 22924 3056 22936
rect 3108 22924 3114 22976
rect 3528 22973 3556 23004
rect 4065 23001 4077 23004
rect 4111 23001 4123 23035
rect 7282 23032 7288 23044
rect 4065 22995 4123 23001
rect 4816 23004 7288 23032
rect 3513 22967 3571 22973
rect 3513 22933 3525 22967
rect 3559 22933 3571 22967
rect 3513 22927 3571 22933
rect 3697 22967 3755 22973
rect 3697 22933 3709 22967
rect 3743 22964 3755 22967
rect 4816 22964 4844 23004
rect 7282 22992 7288 23004
rect 7340 22992 7346 23044
rect 21450 23032 21456 23044
rect 16684 23004 21456 23032
rect 16684 22976 16712 23004
rect 21450 22992 21456 23004
rect 21508 22992 21514 23044
rect 3743 22936 4844 22964
rect 3743 22933 3755 22936
rect 3697 22927 3755 22933
rect 7190 22924 7196 22976
rect 7248 22964 7254 22976
rect 9582 22964 9588 22976
rect 7248 22936 9588 22964
rect 7248 22924 7254 22936
rect 9582 22924 9588 22936
rect 9640 22964 9646 22976
rect 11333 22967 11391 22973
rect 11333 22964 11345 22967
rect 9640 22936 11345 22964
rect 9640 22924 9646 22936
rect 11333 22933 11345 22936
rect 11379 22964 11391 22967
rect 14090 22964 14096 22976
rect 11379 22936 14096 22964
rect 11379 22933 11391 22936
rect 11333 22927 11391 22933
rect 14090 22924 14096 22936
rect 14148 22924 14154 22976
rect 16666 22924 16672 22976
rect 16724 22924 16730 22976
rect 18322 22924 18328 22976
rect 18380 22924 18386 22976
rect 552 22874 23368 22896
rect 552 22822 3662 22874
rect 3714 22822 3726 22874
rect 3778 22822 3790 22874
rect 3842 22822 3854 22874
rect 3906 22822 3918 22874
rect 3970 22822 23368 22874
rect 552 22800 23368 22822
rect 4706 22720 4712 22772
rect 4764 22760 4770 22772
rect 7190 22760 7196 22772
rect 4764 22732 7196 22760
rect 4764 22720 4770 22732
rect 7190 22720 7196 22732
rect 7248 22720 7254 22772
rect 7282 22720 7288 22772
rect 7340 22760 7346 22772
rect 7653 22763 7711 22769
rect 7653 22760 7665 22763
rect 7340 22732 7665 22760
rect 7340 22720 7346 22732
rect 7653 22729 7665 22732
rect 7699 22760 7711 22763
rect 8202 22760 8208 22772
rect 7699 22732 8208 22760
rect 7699 22729 7711 22732
rect 7653 22723 7711 22729
rect 8202 22720 8208 22732
rect 8260 22720 8266 22772
rect 12069 22763 12127 22769
rect 10428 22732 11836 22760
rect 5994 22692 6000 22704
rect 3804 22664 6000 22692
rect 3804 22633 3832 22664
rect 5994 22652 6000 22664
rect 6052 22652 6058 22704
rect 10428 22692 10456 22732
rect 7852 22664 10456 22692
rect 10505 22695 10563 22701
rect 3789 22627 3847 22633
rect 3068 22596 3648 22624
rect 3068 22568 3096 22596
rect 3050 22516 3056 22568
rect 3108 22516 3114 22568
rect 3418 22516 3424 22568
rect 3476 22516 3482 22568
rect 3620 22565 3648 22596
rect 3789 22593 3801 22627
rect 3835 22593 3847 22627
rect 3789 22587 3847 22593
rect 7852 22568 7880 22664
rect 10505 22661 10517 22695
rect 10551 22661 10563 22695
rect 11808 22692 11836 22732
rect 12069 22729 12081 22763
rect 12115 22760 12127 22763
rect 12621 22763 12679 22769
rect 12621 22760 12633 22763
rect 12115 22732 12633 22760
rect 12115 22729 12127 22732
rect 12069 22723 12127 22729
rect 12621 22729 12633 22732
rect 12667 22760 12679 22763
rect 13998 22760 14004 22772
rect 12667 22732 14004 22760
rect 12667 22729 12679 22732
rect 12621 22723 12679 22729
rect 13998 22720 14004 22732
rect 14056 22720 14062 22772
rect 15286 22720 15292 22772
rect 15344 22760 15350 22772
rect 17589 22763 17647 22769
rect 15344 22732 15976 22760
rect 15344 22720 15350 22732
rect 15197 22695 15255 22701
rect 11808 22664 13952 22692
rect 10505 22655 10563 22661
rect 10520 22624 10548 22655
rect 13814 22624 13820 22636
rect 10520 22596 13820 22624
rect 3605 22559 3663 22565
rect 3605 22525 3617 22559
rect 3651 22525 3663 22559
rect 3605 22519 3663 22525
rect 4065 22559 4123 22565
rect 4065 22525 4077 22559
rect 4111 22556 4123 22559
rect 4338 22556 4344 22568
rect 4111 22528 4344 22556
rect 4111 22525 4123 22528
rect 4065 22519 4123 22525
rect 4338 22516 4344 22528
rect 4396 22516 4402 22568
rect 4706 22516 4712 22568
rect 4764 22516 4770 22568
rect 4798 22516 4804 22568
rect 4856 22556 4862 22568
rect 5000 22565 5212 22566
rect 5000 22559 5227 22565
rect 5000 22556 5181 22559
rect 4856 22538 5181 22556
rect 4856 22528 5028 22538
rect 4856 22516 4862 22528
rect 5169 22525 5181 22538
rect 5215 22525 5227 22559
rect 5169 22519 5227 22525
rect 6270 22516 6276 22568
rect 6328 22556 6334 22568
rect 7285 22559 7343 22565
rect 7285 22556 7297 22559
rect 6328 22528 7297 22556
rect 6328 22516 6334 22528
rect 7285 22525 7297 22528
rect 7331 22556 7343 22559
rect 7466 22556 7472 22568
rect 7331 22528 7472 22556
rect 7331 22525 7343 22528
rect 7285 22519 7343 22525
rect 7466 22516 7472 22528
rect 7524 22516 7530 22568
rect 7653 22559 7711 22565
rect 7653 22525 7665 22559
rect 7699 22556 7711 22559
rect 7834 22556 7840 22568
rect 7699 22528 7840 22556
rect 7699 22525 7711 22528
rect 7653 22519 7711 22525
rect 7834 22516 7840 22528
rect 7892 22516 7898 22568
rect 8478 22516 8484 22568
rect 8536 22556 8542 22568
rect 8757 22559 8815 22565
rect 8757 22556 8769 22559
rect 8536 22528 8769 22556
rect 8536 22516 8542 22528
rect 8757 22525 8769 22528
rect 8803 22525 8815 22559
rect 8757 22519 8815 22525
rect 10229 22559 10287 22565
rect 10229 22525 10241 22559
rect 10275 22556 10287 22559
rect 10594 22556 10600 22568
rect 10275 22528 10600 22556
rect 10275 22525 10287 22528
rect 10229 22519 10287 22525
rect 10594 22516 10600 22528
rect 10652 22516 10658 22568
rect 11790 22516 11796 22568
rect 11848 22516 11854 22568
rect 12526 22516 12532 22568
rect 12584 22516 12590 22568
rect 12636 22565 12664 22596
rect 13814 22584 13820 22596
rect 13872 22584 13878 22636
rect 12621 22559 12679 22565
rect 12621 22525 12633 22559
rect 12667 22525 12679 22559
rect 12621 22519 12679 22525
rect 12713 22559 12771 22565
rect 12713 22525 12725 22559
rect 12759 22525 12771 22559
rect 12713 22519 12771 22525
rect 5080 22500 5132 22506
rect 7742 22448 7748 22500
rect 7800 22488 7806 22500
rect 8389 22491 8447 22497
rect 8389 22488 8401 22491
rect 7800 22460 8401 22488
rect 7800 22448 7806 22460
rect 8389 22457 8401 22460
rect 8435 22457 8447 22491
rect 8389 22451 8447 22457
rect 8573 22491 8631 22497
rect 8573 22457 8585 22491
rect 8619 22457 8631 22491
rect 8573 22451 8631 22457
rect 5080 22442 5132 22448
rect 2866 22380 2872 22432
rect 2924 22380 2930 22432
rect 7098 22380 7104 22432
rect 7156 22420 7162 22432
rect 7469 22423 7527 22429
rect 7469 22420 7481 22423
rect 7156 22392 7481 22420
rect 7156 22380 7162 22392
rect 7469 22389 7481 22392
rect 7515 22420 7527 22423
rect 7926 22420 7932 22432
rect 7515 22392 7932 22420
rect 7515 22389 7527 22392
rect 7469 22383 7527 22389
rect 7926 22380 7932 22392
rect 7984 22380 7990 22432
rect 8202 22380 8208 22432
rect 8260 22420 8266 22432
rect 8588 22420 8616 22451
rect 10410 22448 10416 22500
rect 10468 22488 10474 22500
rect 10505 22491 10563 22497
rect 10505 22488 10517 22491
rect 10468 22460 10517 22488
rect 10468 22448 10474 22460
rect 10505 22457 10517 22460
rect 10551 22457 10563 22491
rect 10505 22451 10563 22457
rect 12066 22448 12072 22500
rect 12124 22448 12130 22500
rect 12434 22448 12440 22500
rect 12492 22488 12498 22500
rect 12728 22488 12756 22519
rect 12802 22516 12808 22568
rect 12860 22516 12866 22568
rect 12894 22488 12900 22500
rect 12492 22460 12900 22488
rect 12492 22448 12498 22460
rect 12894 22448 12900 22460
rect 12952 22448 12958 22500
rect 8662 22420 8668 22432
rect 8260 22392 8668 22420
rect 8260 22380 8266 22392
rect 8662 22380 8668 22392
rect 8720 22380 8726 22432
rect 10318 22380 10324 22432
rect 10376 22380 10382 22432
rect 11698 22380 11704 22432
rect 11756 22420 11762 22432
rect 11885 22423 11943 22429
rect 11885 22420 11897 22423
rect 11756 22392 11897 22420
rect 11756 22380 11762 22392
rect 11885 22389 11897 22392
rect 11931 22389 11943 22423
rect 11885 22383 11943 22389
rect 12250 22380 12256 22432
rect 12308 22380 12314 22432
rect 12710 22380 12716 22432
rect 12768 22420 12774 22432
rect 13081 22423 13139 22429
rect 13081 22420 13093 22423
rect 12768 22392 13093 22420
rect 12768 22380 12774 22392
rect 13081 22389 13093 22392
rect 13127 22389 13139 22423
rect 13081 22383 13139 22389
rect 13725 22423 13783 22429
rect 13725 22389 13737 22423
rect 13771 22420 13783 22423
rect 13924 22420 13952 22664
rect 15197 22661 15209 22695
rect 15243 22692 15255 22695
rect 15948 22692 15976 22732
rect 17589 22729 17601 22763
rect 17635 22729 17647 22763
rect 17589 22723 17647 22729
rect 17773 22763 17831 22769
rect 17773 22729 17785 22763
rect 17819 22760 17831 22763
rect 17954 22760 17960 22772
rect 17819 22732 17960 22760
rect 17819 22729 17831 22732
rect 17773 22723 17831 22729
rect 17604 22692 17632 22723
rect 17954 22720 17960 22732
rect 18012 22720 18018 22772
rect 20625 22695 20683 22701
rect 15243 22664 15516 22692
rect 15243 22661 15255 22664
rect 15197 22655 15255 22661
rect 14001 22627 14059 22633
rect 14001 22593 14013 22627
rect 14047 22593 14059 22627
rect 14001 22587 14059 22593
rect 14108 22596 15424 22624
rect 14016 22488 14044 22587
rect 14108 22568 14136 22596
rect 14090 22516 14096 22568
rect 14148 22516 14154 22568
rect 14921 22559 14979 22565
rect 14921 22525 14933 22559
rect 14967 22556 14979 22559
rect 15286 22556 15292 22568
rect 14967 22528 15292 22556
rect 14967 22525 14979 22528
rect 14921 22519 14979 22525
rect 14182 22488 14188 22500
rect 14016 22460 14188 22488
rect 14182 22448 14188 22460
rect 14240 22488 14246 22500
rect 14936 22488 14964 22519
rect 15286 22516 15292 22528
rect 15344 22516 15350 22568
rect 14240 22460 14964 22488
rect 14240 22448 14246 22460
rect 15194 22448 15200 22500
rect 15252 22448 15258 22500
rect 14826 22420 14832 22432
rect 13771 22392 14832 22420
rect 13771 22389 13783 22392
rect 13725 22383 13783 22389
rect 14826 22380 14832 22392
rect 14884 22380 14890 22432
rect 15010 22380 15016 22432
rect 15068 22380 15074 22432
rect 15286 22380 15292 22432
rect 15344 22380 15350 22432
rect 15396 22420 15424 22596
rect 15488 22565 15516 22664
rect 15948 22664 20484 22692
rect 15948 22633 15976 22664
rect 15933 22627 15991 22633
rect 15933 22593 15945 22627
rect 15979 22593 15991 22627
rect 15933 22587 15991 22593
rect 15473 22559 15531 22565
rect 15473 22525 15485 22559
rect 15519 22556 15531 22559
rect 16850 22556 16856 22568
rect 15519 22528 16856 22556
rect 15519 22525 15531 22528
rect 15473 22519 15531 22525
rect 16850 22516 16856 22528
rect 16908 22516 16914 22568
rect 17880 22565 17908 22664
rect 18322 22584 18328 22636
rect 18380 22624 18386 22636
rect 18877 22627 18935 22633
rect 18877 22624 18889 22627
rect 18380 22596 18889 22624
rect 18380 22584 18386 22596
rect 18877 22593 18889 22596
rect 18923 22593 18935 22627
rect 18877 22587 18935 22593
rect 17865 22559 17923 22565
rect 17865 22525 17877 22559
rect 17911 22525 17923 22559
rect 17865 22519 17923 22525
rect 18049 22559 18107 22565
rect 18049 22525 18061 22559
rect 18095 22525 18107 22559
rect 18414 22556 18420 22568
rect 18049 22519 18107 22525
rect 18156 22528 18420 22556
rect 15654 22448 15660 22500
rect 15712 22448 15718 22500
rect 16666 22448 16672 22500
rect 16724 22448 16730 22500
rect 17405 22491 17463 22497
rect 17405 22457 17417 22491
rect 17451 22488 17463 22491
rect 18064 22488 18092 22519
rect 17451 22460 18092 22488
rect 17451 22457 17463 22460
rect 17405 22451 17463 22457
rect 17420 22420 17448 22451
rect 15396 22392 17448 22420
rect 17615 22423 17673 22429
rect 17615 22389 17627 22423
rect 17661 22420 17673 22423
rect 18156 22420 18184 22528
rect 18414 22516 18420 22528
rect 18472 22516 18478 22568
rect 18969 22559 19027 22565
rect 18969 22525 18981 22559
rect 19015 22556 19027 22559
rect 19242 22556 19248 22568
rect 19015 22528 19248 22556
rect 19015 22525 19027 22528
rect 18969 22519 19027 22525
rect 19242 22516 19248 22528
rect 19300 22516 19306 22568
rect 19797 22559 19855 22565
rect 19797 22525 19809 22559
rect 19843 22556 19855 22559
rect 20070 22556 20076 22568
rect 19843 22528 20076 22556
rect 19843 22525 19855 22528
rect 19797 22519 19855 22525
rect 20070 22516 20076 22528
rect 20128 22556 20134 22568
rect 20349 22559 20407 22565
rect 20349 22556 20361 22559
rect 20128 22528 20361 22556
rect 20128 22516 20134 22528
rect 20349 22525 20361 22528
rect 20395 22525 20407 22559
rect 20456 22556 20484 22664
rect 20625 22661 20637 22695
rect 20671 22692 20683 22695
rect 20671 22664 21772 22692
rect 20671 22661 20683 22664
rect 20625 22655 20683 22661
rect 20714 22584 20720 22636
rect 20772 22624 20778 22636
rect 20901 22627 20959 22633
rect 20901 22624 20913 22627
rect 20772 22596 20913 22624
rect 20772 22584 20778 22596
rect 20901 22593 20913 22596
rect 20947 22593 20959 22627
rect 20901 22587 20959 22593
rect 21358 22584 21364 22636
rect 21416 22584 21422 22636
rect 21744 22565 21772 22664
rect 21269 22559 21327 22565
rect 21269 22556 21281 22559
rect 20456 22528 21281 22556
rect 20349 22519 20407 22525
rect 21269 22525 21281 22528
rect 21315 22525 21327 22559
rect 21269 22519 21327 22525
rect 21729 22559 21787 22565
rect 21729 22525 21741 22559
rect 21775 22525 21787 22559
rect 21729 22519 21787 22525
rect 20622 22448 20628 22500
rect 20680 22448 20686 22500
rect 20806 22448 20812 22500
rect 20864 22488 20870 22500
rect 21818 22488 21824 22500
rect 20864 22460 21824 22488
rect 20864 22448 20870 22460
rect 21818 22448 21824 22460
rect 21876 22488 21882 22500
rect 21913 22491 21971 22497
rect 21913 22488 21925 22491
rect 21876 22460 21925 22488
rect 21876 22448 21882 22460
rect 21913 22457 21925 22460
rect 21959 22457 21971 22491
rect 21913 22451 21971 22457
rect 17661 22392 18184 22420
rect 18325 22423 18383 22429
rect 17661 22389 17673 22392
rect 17615 22383 17673 22389
rect 18325 22389 18337 22423
rect 18371 22420 18383 22423
rect 18782 22420 18788 22432
rect 18371 22392 18788 22420
rect 18371 22389 18383 22392
rect 18325 22383 18383 22389
rect 18782 22380 18788 22392
rect 18840 22380 18846 22432
rect 19886 22380 19892 22432
rect 19944 22420 19950 22432
rect 20441 22423 20499 22429
rect 20441 22420 20453 22423
rect 19944 22392 20453 22420
rect 19944 22380 19950 22392
rect 20441 22389 20453 22392
rect 20487 22389 20499 22423
rect 20441 22383 20499 22389
rect 21542 22380 21548 22432
rect 21600 22380 21606 22432
rect 552 22330 23368 22352
rect 552 22278 4322 22330
rect 4374 22278 4386 22330
rect 4438 22278 4450 22330
rect 4502 22278 4514 22330
rect 4566 22278 4578 22330
rect 4630 22278 23368 22330
rect 552 22256 23368 22278
rect 6822 22216 6828 22228
rect 6656 22188 6828 22216
rect 6270 22148 6276 22160
rect 5828 22120 6276 22148
rect 5828 22092 5856 22120
rect 6270 22108 6276 22120
rect 6328 22108 6334 22160
rect 6473 22151 6531 22157
rect 6473 22148 6485 22151
rect 6380 22120 6485 22148
rect 4246 22040 4252 22092
rect 4304 22040 4310 22092
rect 5074 22040 5080 22092
rect 5132 22040 5138 22092
rect 5810 22040 5816 22092
rect 5868 22040 5874 22092
rect 5994 22040 6000 22092
rect 6052 22080 6058 22092
rect 6380 22080 6408 22120
rect 6473 22117 6485 22120
rect 6519 22148 6531 22151
rect 6656 22148 6684 22188
rect 6822 22176 6828 22188
rect 6880 22176 6886 22228
rect 8478 22176 8484 22228
rect 8536 22176 8542 22228
rect 12526 22176 12532 22228
rect 12584 22216 12590 22228
rect 13354 22216 13360 22228
rect 12584 22188 13360 22216
rect 12584 22176 12590 22188
rect 13354 22176 13360 22188
rect 13412 22176 13418 22228
rect 13906 22176 13912 22228
rect 13964 22216 13970 22228
rect 14090 22216 14096 22228
rect 13964 22188 14096 22216
rect 13964 22176 13970 22188
rect 14090 22176 14096 22188
rect 14148 22216 14154 22228
rect 15010 22216 15016 22228
rect 14148 22188 15016 22216
rect 14148 22176 14154 22188
rect 15010 22176 15016 22188
rect 15068 22216 15074 22228
rect 15068 22188 15608 22216
rect 15068 22176 15074 22188
rect 7377 22151 7435 22157
rect 7377 22148 7389 22151
rect 6519 22120 6684 22148
rect 6748 22120 7389 22148
rect 6519 22117 6531 22120
rect 6473 22111 6531 22117
rect 6748 22089 6776 22120
rect 7377 22117 7389 22120
rect 7423 22148 7435 22151
rect 8110 22148 8116 22160
rect 7423 22120 8116 22148
rect 7423 22117 7435 22120
rect 7377 22111 7435 22117
rect 8110 22108 8116 22120
rect 8168 22108 8174 22160
rect 8496 22148 8524 22176
rect 11790 22148 11796 22160
rect 8220 22120 8432 22148
rect 8496 22120 9536 22148
rect 6052 22052 6408 22080
rect 6733 22083 6791 22089
rect 6052 22040 6058 22052
rect 6733 22049 6745 22083
rect 6779 22049 6791 22083
rect 6733 22043 6791 22049
rect 6825 22083 6883 22089
rect 6825 22049 6837 22083
rect 6871 22049 6883 22083
rect 6825 22043 6883 22049
rect 6840 22012 6868 22043
rect 7006 22040 7012 22092
rect 7064 22040 7070 22092
rect 7098 22040 7104 22092
rect 7156 22040 7162 22092
rect 7742 22040 7748 22092
rect 7800 22040 7806 22092
rect 7926 22040 7932 22092
rect 7984 22080 7990 22092
rect 8021 22083 8079 22089
rect 8021 22080 8033 22083
rect 7984 22052 8033 22080
rect 7984 22040 7990 22052
rect 8021 22049 8033 22052
rect 8067 22080 8079 22083
rect 8220 22080 8248 22120
rect 8067 22052 8248 22080
rect 8067 22049 8079 22052
rect 8021 22043 8079 22049
rect 8294 22040 8300 22092
rect 8352 22040 8358 22092
rect 8404 22080 8432 22120
rect 9508 22092 9536 22120
rect 10244 22120 11796 22148
rect 8481 22083 8539 22089
rect 8481 22080 8493 22083
rect 8404 22052 8493 22080
rect 8481 22049 8493 22052
rect 8527 22049 8539 22083
rect 8481 22043 8539 22049
rect 8570 22040 8576 22092
rect 8628 22040 8634 22092
rect 8662 22040 8668 22092
rect 8720 22040 8726 22092
rect 9306 22040 9312 22092
rect 9364 22040 9370 22092
rect 9490 22080 9496 22092
rect 9471 22052 9496 22080
rect 9490 22040 9496 22052
rect 9548 22040 9554 22092
rect 6914 22012 6920 22024
rect 6840 21984 6920 22012
rect 5166 21904 5172 21956
rect 5224 21904 5230 21956
rect 6641 21947 6699 21953
rect 6641 21913 6653 21947
rect 6687 21944 6699 21947
rect 6840 21944 6868 21984
rect 6914 21972 6920 21984
rect 6972 21972 6978 22024
rect 7024 22012 7052 22040
rect 8113 22015 8171 22021
rect 7024 21984 7144 22012
rect 6687 21916 6868 21944
rect 7116 21944 7144 21984
rect 8113 21981 8125 22015
rect 8159 22012 8171 22015
rect 10244 22012 10272 22120
rect 11790 22108 11796 22120
rect 11848 22148 11854 22160
rect 13509 22151 13567 22157
rect 13509 22148 13521 22151
rect 11848 22120 13521 22148
rect 11848 22108 11854 22120
rect 13509 22117 13521 22120
rect 13555 22117 13567 22151
rect 13509 22111 13567 22117
rect 13722 22108 13728 22160
rect 13780 22148 13786 22160
rect 14734 22148 14740 22160
rect 13780 22120 14740 22148
rect 13780 22108 13786 22120
rect 14734 22108 14740 22120
rect 14792 22108 14798 22160
rect 15304 22157 15332 22188
rect 15289 22151 15347 22157
rect 15289 22117 15301 22151
rect 15335 22117 15347 22151
rect 15289 22111 15347 22117
rect 15470 22108 15476 22160
rect 15528 22157 15534 22160
rect 15528 22151 15547 22157
rect 15535 22117 15547 22151
rect 15580 22148 15608 22188
rect 15654 22176 15660 22228
rect 15712 22176 15718 22228
rect 16942 22176 16948 22228
rect 17000 22216 17006 22228
rect 20099 22219 20157 22225
rect 17000 22188 19932 22216
rect 17000 22176 17006 22188
rect 16960 22148 16988 22176
rect 19904 22160 19932 22188
rect 20099 22185 20111 22219
rect 20145 22216 20157 22219
rect 20622 22216 20628 22228
rect 20145 22188 20628 22216
rect 20145 22185 20157 22188
rect 20099 22179 20157 22185
rect 20622 22176 20628 22188
rect 20680 22176 20686 22228
rect 21358 22176 21364 22228
rect 21416 22216 21422 22228
rect 22002 22216 22008 22228
rect 21416 22188 22008 22216
rect 21416 22176 21422 22188
rect 22002 22176 22008 22188
rect 22060 22216 22066 22228
rect 22060 22188 22784 22216
rect 22060 22176 22066 22188
rect 19242 22148 19248 22160
rect 15580 22120 16988 22148
rect 17052 22120 19248 22148
rect 15528 22111 15547 22117
rect 15528 22108 15534 22111
rect 10410 22040 10416 22092
rect 10468 22040 10474 22092
rect 10502 22040 10508 22092
rect 10560 22080 10566 22092
rect 10560 22052 10605 22080
rect 10560 22040 10566 22052
rect 10778 22040 10784 22092
rect 10836 22080 10842 22092
rect 11057 22083 11115 22089
rect 11057 22080 11069 22083
rect 10836 22052 11069 22080
rect 10836 22040 10842 22052
rect 11057 22049 11069 22052
rect 11103 22049 11115 22083
rect 12069 22083 12127 22089
rect 11057 22043 11115 22049
rect 8159 21984 10272 22012
rect 10321 22015 10379 22021
rect 8159 21981 8171 21984
rect 8113 21975 8171 21981
rect 10321 21981 10333 22015
rect 10367 22012 10379 22015
rect 10686 22012 10692 22024
rect 10367 21984 10692 22012
rect 10367 21981 10379 21984
rect 10321 21975 10379 21981
rect 10686 21972 10692 21984
rect 10744 22012 10750 22024
rect 11164 22012 11192 22066
rect 12069 22049 12081 22083
rect 12115 22080 12127 22083
rect 12529 22083 12587 22089
rect 12529 22080 12541 22083
rect 12115 22052 12541 22080
rect 12115 22049 12127 22052
rect 12069 22043 12127 22049
rect 12529 22049 12541 22052
rect 12575 22080 12587 22083
rect 12802 22080 12808 22092
rect 12575 22052 12808 22080
rect 12575 22049 12587 22052
rect 12529 22043 12587 22049
rect 12802 22040 12808 22052
rect 12860 22040 12866 22092
rect 12894 22040 12900 22092
rect 12952 22040 12958 22092
rect 13354 22040 13360 22092
rect 13412 22080 13418 22092
rect 13412 22052 13952 22080
rect 13412 22040 13418 22052
rect 10744 21984 11192 22012
rect 10744 21972 10750 21984
rect 13262 21972 13268 22024
rect 13320 21972 13326 22024
rect 13814 21972 13820 22024
rect 13872 21972 13878 22024
rect 13924 22012 13952 22052
rect 13998 22040 14004 22092
rect 14056 22040 14062 22092
rect 14093 22083 14151 22089
rect 14093 22049 14105 22083
rect 14139 22049 14151 22083
rect 14093 22043 14151 22049
rect 15013 22083 15071 22089
rect 15013 22049 15025 22083
rect 15059 22049 15071 22083
rect 15013 22043 15071 22049
rect 14108 22012 14136 22043
rect 13924 21984 14136 22012
rect 15028 21956 15056 22043
rect 15654 22040 15660 22092
rect 15712 22080 15718 22092
rect 16117 22083 16175 22089
rect 16117 22080 16129 22083
rect 15712 22052 16129 22080
rect 15712 22040 15718 22052
rect 16117 22049 16129 22052
rect 16163 22049 16175 22083
rect 16117 22043 16175 22049
rect 16850 22040 16856 22092
rect 16908 22040 16914 22092
rect 17052 22089 17080 22120
rect 19242 22108 19248 22120
rect 19300 22108 19306 22160
rect 19886 22108 19892 22160
rect 19944 22108 19950 22160
rect 21376 22148 21404 22176
rect 22756 22157 22784 22188
rect 22557 22151 22615 22157
rect 22557 22148 22569 22151
rect 20824 22120 21404 22148
rect 22020 22126 22569 22148
rect 17037 22083 17095 22089
rect 17037 22049 17049 22083
rect 17083 22049 17095 22083
rect 17037 22043 17095 22049
rect 17681 22083 17739 22089
rect 17681 22049 17693 22083
rect 17727 22049 17739 22083
rect 17681 22043 17739 22049
rect 15105 22015 15163 22021
rect 15105 21981 15117 22015
rect 15151 22012 15163 22015
rect 15286 22012 15292 22024
rect 15151 21984 15292 22012
rect 15151 21981 15163 21984
rect 15105 21975 15163 21981
rect 15286 21972 15292 21984
rect 15344 21972 15350 22024
rect 16666 21972 16672 22024
rect 16724 22012 16730 22024
rect 17052 22012 17080 22043
rect 16724 21984 17080 22012
rect 17696 22012 17724 22043
rect 17954 22040 17960 22092
rect 18012 22080 18018 22092
rect 18141 22083 18199 22089
rect 18141 22080 18153 22083
rect 18012 22052 18153 22080
rect 18012 22040 18018 22052
rect 18141 22049 18153 22052
rect 18187 22049 18199 22083
rect 18141 22043 18199 22049
rect 18782 22040 18788 22092
rect 18840 22040 18846 22092
rect 20824 22080 20852 22120
rect 20456 22052 20852 22080
rect 20901 22083 20959 22089
rect 18046 22012 18052 22024
rect 17696 21984 18052 22012
rect 16724 21972 16730 21984
rect 18046 21972 18052 21984
rect 18104 21972 18110 22024
rect 18322 21972 18328 22024
rect 18380 22012 18386 22024
rect 20346 22012 20352 22024
rect 18380 21984 20352 22012
rect 18380 21972 18386 21984
rect 20346 21972 20352 21984
rect 20404 21972 20410 22024
rect 8205 21947 8263 21953
rect 8205 21944 8217 21947
rect 7116 21916 8217 21944
rect 6687 21913 6699 21916
rect 6641 21907 6699 21913
rect 8205 21913 8217 21916
rect 8251 21913 8263 21947
rect 8205 21907 8263 21913
rect 8941 21947 8999 21953
rect 8941 21913 8953 21947
rect 8987 21944 8999 21947
rect 10410 21944 10416 21956
rect 8987 21916 10416 21944
rect 8987 21913 8999 21916
rect 8941 21907 8999 21913
rect 10410 21904 10416 21916
rect 10468 21904 10474 21956
rect 11698 21904 11704 21956
rect 11756 21944 11762 21956
rect 11756 21916 12940 21944
rect 11756 21904 11762 21916
rect 5902 21836 5908 21888
rect 5960 21836 5966 21888
rect 6362 21836 6368 21888
rect 6420 21876 6426 21888
rect 6457 21879 6515 21885
rect 6457 21876 6469 21879
rect 6420 21848 6469 21876
rect 6420 21836 6426 21848
rect 6457 21845 6469 21848
rect 6503 21845 6515 21879
rect 6457 21839 6515 21845
rect 7282 21836 7288 21888
rect 7340 21836 7346 21888
rect 10226 21836 10232 21888
rect 10284 21876 10290 21888
rect 10597 21879 10655 21885
rect 10597 21876 10609 21879
rect 10284 21848 10609 21876
rect 10284 21836 10290 21848
rect 10597 21845 10609 21848
rect 10643 21845 10655 21879
rect 12912 21876 12940 21916
rect 14642 21904 14648 21956
rect 14700 21904 14706 21956
rect 15010 21904 15016 21956
rect 15068 21944 15074 21956
rect 20456 21944 20484 22052
rect 20901 22049 20913 22083
rect 20947 22049 20959 22083
rect 20901 22043 20959 22049
rect 21085 22083 21143 22089
rect 21085 22049 21097 22083
rect 21131 22049 21143 22083
rect 21376 22080 21404 22120
rect 21634 22080 21640 22092
rect 21376 22052 21640 22080
rect 21085 22043 21143 22049
rect 20809 22015 20867 22021
rect 20809 21981 20821 22015
rect 20855 22012 20867 22015
rect 20916 22012 20944 22043
rect 20855 21984 20944 22012
rect 20855 21981 20867 21984
rect 20809 21975 20867 21981
rect 21100 21956 21128 22043
rect 21634 22040 21640 22052
rect 21692 22040 21698 22092
rect 21818 22040 21824 22092
rect 21876 22080 21882 22092
rect 21913 22083 21971 22089
rect 21913 22080 21925 22083
rect 21876 22052 21925 22080
rect 21876 22040 21882 22052
rect 21913 22049 21925 22052
rect 21959 22049 21971 22083
rect 22002 22074 22008 22126
rect 22060 22120 22569 22126
rect 22060 22074 22066 22120
rect 22557 22117 22569 22120
rect 22603 22117 22615 22151
rect 22557 22111 22615 22117
rect 22741 22151 22799 22157
rect 22741 22117 22753 22151
rect 22787 22117 22799 22151
rect 22741 22111 22799 22117
rect 21913 22043 21971 22049
rect 22094 22040 22100 22092
rect 22152 22080 22158 22092
rect 22465 22083 22523 22089
rect 22465 22080 22477 22083
rect 22152 22052 22477 22080
rect 22152 22040 22158 22052
rect 22465 22049 22477 22052
rect 22511 22049 22523 22083
rect 22465 22043 22523 22049
rect 21450 21972 21456 22024
rect 21508 22012 21514 22024
rect 22002 22012 22008 22024
rect 21508 21984 22008 22012
rect 21508 21972 21514 21984
rect 22002 21972 22008 21984
rect 22060 21972 22066 22024
rect 22189 22015 22247 22021
rect 22189 21981 22201 22015
rect 22235 21981 22247 22015
rect 22189 21975 22247 21981
rect 15068 21916 20484 21944
rect 20625 21947 20683 21953
rect 15068 21904 15074 21916
rect 20625 21913 20637 21947
rect 20671 21944 20683 21947
rect 20714 21944 20720 21956
rect 20671 21916 20720 21944
rect 20671 21913 20683 21916
rect 20625 21907 20683 21913
rect 20714 21904 20720 21916
rect 20772 21944 20778 21956
rect 20990 21944 20996 21956
rect 20772 21916 20996 21944
rect 20772 21904 20778 21916
rect 20990 21904 20996 21916
rect 21048 21904 21054 21956
rect 21082 21904 21088 21956
rect 21140 21944 21146 21956
rect 21140 21916 21496 21944
rect 21140 21904 21146 21916
rect 13541 21879 13599 21885
rect 13541 21876 13553 21879
rect 12912 21848 13553 21876
rect 10597 21839 10655 21845
rect 13541 21845 13553 21848
rect 13587 21845 13599 21879
rect 13541 21839 13599 21845
rect 13722 21836 13728 21888
rect 13780 21876 13786 21888
rect 13909 21879 13967 21885
rect 13909 21876 13921 21879
rect 13780 21848 13921 21876
rect 13780 21836 13786 21848
rect 13909 21845 13921 21848
rect 13955 21845 13967 21879
rect 13909 21839 13967 21845
rect 14182 21836 14188 21888
rect 14240 21876 14246 21888
rect 15473 21879 15531 21885
rect 15473 21876 15485 21879
rect 14240 21848 15485 21876
rect 14240 21836 14246 21848
rect 15473 21845 15485 21848
rect 15519 21845 15531 21879
rect 15473 21839 15531 21845
rect 16298 21836 16304 21888
rect 16356 21836 16362 21888
rect 17773 21879 17831 21885
rect 17773 21845 17785 21879
rect 17819 21876 17831 21879
rect 18138 21876 18144 21888
rect 17819 21848 18144 21876
rect 17819 21845 17831 21848
rect 17773 21839 17831 21845
rect 18138 21836 18144 21848
rect 18196 21836 18202 21888
rect 18322 21836 18328 21888
rect 18380 21836 18386 21888
rect 19242 21836 19248 21888
rect 19300 21876 19306 21888
rect 19429 21879 19487 21885
rect 19429 21876 19441 21879
rect 19300 21848 19441 21876
rect 19300 21836 19306 21848
rect 19429 21845 19441 21848
rect 19475 21845 19487 21879
rect 19429 21839 19487 21845
rect 19518 21836 19524 21888
rect 19576 21876 19582 21888
rect 20070 21876 20076 21888
rect 19576 21848 20076 21876
rect 19576 21836 19582 21848
rect 20070 21836 20076 21848
rect 20128 21836 20134 21888
rect 20257 21879 20315 21885
rect 20257 21845 20269 21879
rect 20303 21876 20315 21879
rect 20806 21876 20812 21888
rect 20303 21848 20812 21876
rect 20303 21845 20315 21848
rect 20257 21839 20315 21845
rect 20806 21836 20812 21848
rect 20864 21836 20870 21888
rect 20898 21836 20904 21888
rect 20956 21836 20962 21888
rect 21174 21836 21180 21888
rect 21232 21876 21238 21888
rect 21361 21879 21419 21885
rect 21361 21876 21373 21879
rect 21232 21848 21373 21876
rect 21232 21836 21238 21848
rect 21361 21845 21373 21848
rect 21407 21845 21419 21879
rect 21468 21876 21496 21916
rect 21726 21904 21732 21956
rect 21784 21944 21790 21956
rect 22204 21944 22232 21975
rect 22278 21972 22284 22024
rect 22336 21972 22342 22024
rect 22465 21947 22523 21953
rect 22465 21944 22477 21947
rect 21784 21916 22477 21944
rect 21784 21904 21790 21916
rect 22465 21913 22477 21916
rect 22511 21913 22523 21947
rect 22465 21907 22523 21913
rect 22005 21879 22063 21885
rect 22005 21876 22017 21879
rect 21468 21848 22017 21876
rect 21361 21839 21419 21845
rect 22005 21845 22017 21848
rect 22051 21845 22063 21879
rect 22005 21839 22063 21845
rect 22094 21836 22100 21888
rect 22152 21836 22158 21888
rect 552 21786 23368 21808
rect 552 21734 3662 21786
rect 3714 21734 3726 21786
rect 3778 21734 3790 21786
rect 3842 21734 3854 21786
rect 3906 21734 3918 21786
rect 3970 21734 23368 21786
rect 552 21712 23368 21734
rect 6914 21632 6920 21684
rect 6972 21672 6978 21684
rect 7742 21672 7748 21684
rect 6972 21644 7748 21672
rect 6972 21632 6978 21644
rect 7742 21632 7748 21644
rect 7800 21632 7806 21684
rect 8110 21632 8116 21684
rect 8168 21672 8174 21684
rect 8205 21675 8263 21681
rect 8205 21672 8217 21675
rect 8168 21644 8217 21672
rect 8168 21632 8174 21644
rect 8205 21641 8217 21644
rect 8251 21672 8263 21675
rect 8570 21672 8576 21684
rect 8251 21644 8576 21672
rect 8251 21641 8263 21644
rect 8205 21635 8263 21641
rect 8570 21632 8576 21644
rect 8628 21632 8634 21684
rect 9766 21632 9772 21684
rect 9824 21672 9830 21684
rect 10502 21672 10508 21684
rect 9824 21644 10508 21672
rect 9824 21632 9830 21644
rect 10502 21632 10508 21644
rect 10560 21632 10566 21684
rect 11885 21675 11943 21681
rect 11885 21641 11897 21675
rect 11931 21672 11943 21675
rect 12434 21672 12440 21684
rect 11931 21644 12440 21672
rect 11931 21641 11943 21644
rect 11885 21635 11943 21641
rect 12434 21632 12440 21644
rect 12492 21632 12498 21684
rect 12894 21632 12900 21684
rect 12952 21672 12958 21684
rect 13630 21672 13636 21684
rect 12952 21644 13636 21672
rect 12952 21632 12958 21644
rect 13630 21632 13636 21644
rect 13688 21632 13694 21684
rect 14734 21632 14740 21684
rect 14792 21672 14798 21684
rect 15562 21672 15568 21684
rect 14792 21644 15568 21672
rect 14792 21632 14798 21644
rect 15562 21632 15568 21644
rect 15620 21632 15626 21684
rect 16393 21675 16451 21681
rect 16393 21641 16405 21675
rect 16439 21672 16451 21675
rect 16758 21672 16764 21684
rect 16439 21644 16764 21672
rect 16439 21641 16451 21644
rect 16393 21635 16451 21641
rect 16758 21632 16764 21644
rect 16816 21672 16822 21684
rect 17405 21675 17463 21681
rect 17405 21672 17417 21675
rect 16816 21644 17417 21672
rect 16816 21632 16822 21644
rect 17405 21641 17417 21644
rect 17451 21641 17463 21675
rect 17405 21635 17463 21641
rect 20806 21632 20812 21684
rect 20864 21672 20870 21684
rect 21177 21675 21235 21681
rect 21177 21672 21189 21675
rect 20864 21644 21189 21672
rect 20864 21632 20870 21644
rect 21177 21641 21189 21644
rect 21223 21641 21235 21675
rect 21177 21635 21235 21641
rect 21358 21632 21364 21684
rect 21416 21672 21422 21684
rect 21726 21672 21732 21684
rect 21416 21644 21732 21672
rect 21416 21632 21422 21644
rect 21726 21632 21732 21644
rect 21784 21632 21790 21684
rect 22005 21675 22063 21681
rect 22005 21641 22017 21675
rect 22051 21672 22063 21675
rect 22278 21672 22284 21684
rect 22051 21644 22284 21672
rect 22051 21641 22063 21644
rect 22005 21635 22063 21641
rect 7193 21607 7251 21613
rect 7193 21573 7205 21607
rect 7239 21604 7251 21607
rect 7558 21604 7564 21616
rect 7239 21576 7564 21604
rect 7239 21573 7251 21576
rect 7193 21567 7251 21573
rect 7558 21564 7564 21576
rect 7616 21604 7622 21616
rect 8294 21604 8300 21616
rect 7616 21576 8300 21604
rect 7616 21564 7622 21576
rect 8294 21564 8300 21576
rect 8352 21564 8358 21616
rect 8846 21604 8852 21616
rect 8588 21576 8852 21604
rect 5166 21496 5172 21548
rect 5224 21496 5230 21548
rect 6270 21496 6276 21548
rect 6328 21536 6334 21548
rect 6549 21539 6607 21545
rect 6549 21536 6561 21539
rect 6328 21508 6561 21536
rect 6328 21496 6334 21508
rect 6549 21505 6561 21508
rect 6595 21505 6607 21539
rect 6549 21499 6607 21505
rect 6822 21496 6828 21548
rect 6880 21536 6886 21548
rect 7377 21539 7435 21545
rect 7377 21536 7389 21539
rect 6880 21508 7389 21536
rect 6880 21496 6886 21508
rect 7377 21505 7389 21508
rect 7423 21536 7435 21539
rect 7423 21508 7788 21536
rect 7423 21505 7435 21508
rect 7377 21499 7435 21505
rect 4246 21428 4252 21480
rect 4304 21428 4310 21480
rect 4617 21471 4675 21477
rect 4617 21437 4629 21471
rect 4663 21468 4675 21471
rect 4798 21468 4804 21480
rect 4663 21440 4804 21468
rect 4663 21437 4675 21440
rect 4617 21431 4675 21437
rect 4798 21428 4804 21440
rect 4856 21428 4862 21480
rect 5261 21471 5319 21477
rect 5261 21437 5273 21471
rect 5307 21468 5319 21471
rect 5902 21468 5908 21480
rect 5307 21440 5908 21468
rect 5307 21437 5319 21440
rect 5261 21431 5319 21437
rect 5902 21428 5908 21440
rect 5960 21428 5966 21480
rect 7009 21471 7067 21477
rect 7009 21470 7021 21471
rect 6932 21442 7021 21470
rect 3881 21403 3939 21409
rect 3881 21369 3893 21403
rect 3927 21369 3939 21403
rect 4816 21400 4844 21428
rect 6932 21400 6960 21442
rect 7009 21437 7021 21442
rect 7055 21437 7067 21471
rect 7009 21431 7067 21437
rect 7024 21406 7060 21431
rect 7466 21428 7472 21480
rect 7524 21468 7530 21480
rect 7650 21468 7656 21480
rect 7524 21440 7656 21468
rect 7524 21428 7530 21440
rect 7650 21428 7656 21440
rect 7708 21428 7714 21480
rect 7760 21468 7788 21508
rect 7834 21496 7840 21548
rect 7892 21496 7898 21548
rect 8588 21536 8616 21576
rect 8846 21564 8852 21576
rect 8904 21564 8910 21616
rect 9490 21564 9496 21616
rect 9548 21604 9554 21616
rect 9677 21607 9735 21613
rect 9677 21604 9689 21607
rect 9548 21576 9689 21604
rect 9548 21564 9554 21576
rect 9677 21573 9689 21576
rect 9723 21573 9735 21607
rect 9677 21567 9735 21573
rect 9861 21607 9919 21613
rect 9861 21573 9873 21607
rect 9907 21604 9919 21607
rect 9907 21576 10916 21604
rect 9907 21573 9919 21576
rect 9861 21567 9919 21573
rect 7944 21508 8616 21536
rect 8680 21508 9168 21536
rect 7944 21477 7972 21508
rect 7929 21471 7987 21477
rect 7929 21468 7941 21471
rect 7760 21440 7941 21468
rect 7929 21437 7941 21440
rect 7975 21437 7987 21471
rect 8128 21468 8340 21470
rect 7929 21431 7987 21437
rect 8036 21442 8524 21468
rect 8036 21440 8156 21442
rect 8312 21440 8524 21442
rect 4816 21372 6960 21400
rect 7032 21400 7060 21406
rect 8036 21400 8064 21440
rect 7032 21372 8064 21400
rect 3881 21363 3939 21369
rect 3896 21332 3924 21363
rect 8202 21360 8208 21412
rect 8260 21400 8266 21412
rect 8496 21400 8524 21440
rect 8570 21428 8576 21480
rect 8628 21428 8634 21480
rect 8680 21400 8708 21508
rect 8846 21428 8852 21480
rect 8904 21428 8910 21480
rect 8938 21428 8944 21480
rect 8996 21428 9002 21480
rect 9140 21477 9168 21508
rect 9214 21496 9220 21548
rect 9272 21536 9278 21548
rect 9309 21539 9367 21545
rect 9309 21536 9321 21539
rect 9272 21508 9321 21536
rect 9272 21496 9278 21508
rect 9309 21505 9321 21508
rect 9355 21536 9367 21539
rect 9582 21536 9588 21548
rect 9355 21508 9588 21536
rect 9355 21505 9367 21508
rect 9309 21499 9367 21505
rect 9582 21496 9588 21508
rect 9640 21496 9646 21548
rect 10226 21496 10232 21548
rect 10284 21496 10290 21548
rect 9125 21471 9183 21477
rect 9125 21437 9137 21471
rect 9171 21462 9183 21471
rect 10137 21471 10195 21477
rect 9171 21437 9260 21462
rect 9125 21434 9260 21437
rect 9125 21431 9183 21434
rect 8260 21372 8305 21400
rect 8496 21372 8708 21400
rect 8757 21403 8815 21409
rect 8260 21360 8266 21372
rect 8757 21369 8769 21403
rect 8803 21400 8815 21403
rect 9030 21400 9036 21412
rect 8803 21372 9036 21400
rect 8803 21369 8815 21372
rect 8757 21363 8815 21369
rect 9030 21360 9036 21372
rect 9088 21360 9094 21412
rect 9232 21400 9260 21434
rect 10137 21437 10149 21471
rect 10183 21468 10195 21471
rect 10318 21468 10324 21480
rect 10183 21440 10324 21468
rect 10183 21437 10195 21440
rect 10137 21431 10195 21437
rect 10318 21428 10324 21440
rect 10376 21428 10382 21480
rect 10597 21471 10655 21477
rect 10597 21437 10609 21471
rect 10643 21468 10655 21471
rect 10686 21468 10692 21480
rect 10643 21440 10692 21468
rect 10643 21437 10655 21440
rect 10597 21431 10655 21437
rect 10686 21428 10692 21440
rect 10744 21428 10750 21480
rect 10888 21477 10916 21576
rect 12526 21564 12532 21616
rect 12584 21604 12590 21616
rect 14090 21604 14096 21616
rect 12584 21576 14096 21604
rect 12584 21564 12590 21576
rect 14090 21564 14096 21576
rect 14148 21564 14154 21616
rect 18322 21604 18328 21616
rect 14660 21576 18328 21604
rect 11698 21496 11704 21548
rect 11756 21496 11762 21548
rect 12250 21496 12256 21548
rect 12308 21496 12314 21548
rect 12710 21496 12716 21548
rect 12768 21496 12774 21548
rect 13722 21536 13728 21548
rect 13004 21508 13728 21536
rect 10873 21471 10931 21477
rect 10873 21437 10885 21471
rect 10919 21437 10931 21471
rect 10873 21431 10931 21437
rect 11790 21428 11796 21480
rect 11848 21468 11854 21480
rect 12161 21471 12219 21477
rect 12161 21468 12173 21471
rect 11848 21440 12173 21468
rect 11848 21428 11854 21440
rect 12161 21437 12173 21440
rect 12207 21437 12219 21471
rect 12161 21431 12219 21437
rect 12437 21471 12495 21477
rect 12437 21437 12449 21471
rect 12483 21470 12495 21471
rect 12483 21468 12664 21470
rect 12802 21468 12808 21480
rect 12483 21442 12808 21468
rect 12483 21437 12495 21442
rect 12636 21440 12808 21442
rect 12437 21431 12495 21437
rect 12802 21428 12808 21440
rect 12860 21468 12866 21480
rect 13004 21468 13032 21508
rect 13722 21496 13728 21508
rect 13780 21496 13786 21548
rect 12860 21440 13032 21468
rect 13081 21471 13139 21477
rect 12860 21428 12866 21440
rect 13081 21437 13093 21471
rect 13127 21437 13139 21471
rect 13081 21431 13139 21437
rect 13173 21471 13231 21477
rect 13173 21437 13185 21471
rect 13219 21468 13231 21471
rect 13262 21468 13268 21480
rect 13219 21440 13268 21468
rect 13219 21437 13231 21440
rect 13173 21431 13231 21437
rect 9306 21400 9312 21412
rect 9232 21372 9312 21400
rect 9306 21360 9312 21372
rect 9364 21360 9370 21412
rect 9398 21360 9404 21412
rect 9456 21360 9462 21412
rect 11330 21400 11336 21412
rect 10520 21372 11336 21400
rect 3970 21332 3976 21344
rect 3896 21304 3976 21332
rect 3970 21292 3976 21304
rect 4028 21292 4034 21344
rect 5902 21292 5908 21344
rect 5960 21292 5966 21344
rect 5997 21335 6055 21341
rect 5997 21301 6009 21335
rect 6043 21332 6055 21335
rect 6178 21332 6184 21344
rect 6043 21304 6184 21332
rect 6043 21301 6055 21304
rect 5997 21295 6055 21301
rect 6178 21292 6184 21304
rect 6236 21292 6242 21344
rect 6362 21292 6368 21344
rect 6420 21292 6426 21344
rect 6457 21335 6515 21341
rect 6457 21301 6469 21335
rect 6503 21332 6515 21335
rect 6917 21335 6975 21341
rect 6917 21332 6929 21335
rect 6503 21304 6929 21332
rect 6503 21301 6515 21304
rect 6457 21295 6515 21301
rect 6917 21301 6929 21304
rect 6963 21301 6975 21335
rect 6917 21295 6975 21301
rect 7742 21292 7748 21344
rect 7800 21332 7806 21344
rect 8021 21335 8079 21341
rect 8021 21332 8033 21335
rect 7800 21304 8033 21332
rect 7800 21292 7806 21304
rect 8021 21301 8033 21304
rect 8067 21301 8079 21335
rect 8021 21295 8079 21301
rect 8389 21335 8447 21341
rect 8389 21301 8401 21335
rect 8435 21332 8447 21335
rect 8570 21332 8576 21344
rect 8435 21304 8576 21332
rect 8435 21301 8447 21304
rect 8389 21295 8447 21301
rect 8570 21292 8576 21304
rect 8628 21292 8634 21344
rect 8662 21292 8668 21344
rect 8720 21332 8726 21344
rect 10134 21332 10140 21344
rect 8720 21304 10140 21332
rect 8720 21292 8726 21304
rect 10134 21292 10140 21304
rect 10192 21292 10198 21344
rect 10520 21341 10548 21372
rect 11330 21360 11336 21372
rect 11388 21360 11394 21412
rect 12066 21360 12072 21412
rect 12124 21400 12130 21412
rect 12894 21400 12900 21412
rect 12124 21372 12900 21400
rect 12124 21360 12130 21372
rect 12894 21360 12900 21372
rect 12952 21360 12958 21412
rect 13096 21400 13124 21431
rect 13262 21428 13268 21440
rect 13320 21468 13326 21480
rect 14553 21471 14611 21477
rect 13320 21440 13938 21468
rect 13320 21428 13326 21440
rect 14553 21437 14565 21471
rect 14599 21468 14611 21471
rect 14660 21468 14688 21576
rect 18322 21564 18328 21576
rect 18380 21564 18386 21616
rect 18417 21607 18475 21613
rect 18417 21573 18429 21607
rect 18463 21604 18475 21607
rect 18463 21576 19564 21604
rect 18463 21573 18475 21576
rect 18417 21567 18475 21573
rect 15289 21539 15347 21545
rect 15289 21536 15301 21539
rect 15028 21508 15301 21536
rect 14599 21440 14688 21468
rect 14599 21437 14611 21440
rect 14553 21431 14611 21437
rect 13096 21372 13492 21400
rect 10505 21335 10563 21341
rect 10505 21301 10517 21335
rect 10551 21301 10563 21335
rect 10505 21295 10563 21301
rect 10686 21292 10692 21344
rect 10744 21292 10750 21344
rect 11054 21292 11060 21344
rect 11112 21292 11118 21344
rect 11146 21292 11152 21344
rect 11204 21332 11210 21344
rect 12526 21332 12532 21344
rect 11204 21304 12532 21332
rect 11204 21292 11210 21304
rect 12526 21292 12532 21304
rect 12584 21292 12590 21344
rect 12621 21335 12679 21341
rect 12621 21301 12633 21335
rect 12667 21332 12679 21335
rect 13078 21332 13084 21344
rect 12667 21304 13084 21332
rect 12667 21301 12679 21304
rect 12621 21295 12679 21301
rect 13078 21292 13084 21304
rect 13136 21292 13142 21344
rect 13354 21292 13360 21344
rect 13412 21292 13418 21344
rect 13464 21332 13492 21372
rect 13538 21360 13544 21412
rect 13596 21360 13602 21412
rect 14660 21332 14688 21440
rect 14826 21428 14832 21480
rect 14884 21468 14890 21480
rect 14921 21471 14979 21477
rect 14921 21468 14933 21471
rect 14884 21440 14933 21468
rect 14884 21428 14890 21440
rect 14921 21437 14933 21440
rect 14967 21437 14979 21471
rect 14921 21431 14979 21437
rect 14734 21360 14740 21412
rect 14792 21360 14798 21412
rect 15028 21400 15056 21508
rect 15289 21505 15301 21508
rect 15335 21505 15347 21539
rect 15289 21499 15347 21505
rect 15562 21496 15568 21548
rect 15620 21536 15626 21548
rect 16853 21539 16911 21545
rect 16853 21536 16865 21539
rect 15620 21508 16865 21536
rect 15620 21496 15626 21508
rect 16853 21505 16865 21508
rect 16899 21536 16911 21539
rect 19426 21536 19432 21548
rect 16899 21508 19432 21536
rect 16899 21505 16911 21508
rect 16853 21499 16911 21505
rect 19426 21496 19432 21508
rect 19484 21496 19490 21548
rect 19536 21480 19564 21576
rect 20346 21564 20352 21616
rect 20404 21604 20410 21616
rect 20717 21607 20775 21613
rect 20717 21604 20729 21607
rect 20404 21576 20729 21604
rect 20404 21564 20410 21576
rect 20717 21573 20729 21576
rect 20763 21573 20775 21607
rect 20717 21567 20775 21573
rect 20901 21607 20959 21613
rect 20901 21573 20913 21607
rect 20947 21573 20959 21607
rect 20901 21567 20959 21573
rect 20916 21536 20944 21567
rect 20990 21564 20996 21616
rect 21048 21604 21054 21616
rect 21542 21604 21548 21616
rect 21048 21576 21548 21604
rect 21048 21564 21054 21576
rect 21542 21564 21548 21576
rect 21600 21564 21606 21616
rect 21082 21536 21088 21548
rect 20916 21508 21088 21536
rect 21082 21496 21088 21508
rect 21140 21496 21146 21548
rect 22020 21536 22048 21635
rect 22278 21632 22284 21644
rect 22336 21632 22342 21684
rect 21468 21508 22048 21536
rect 15102 21428 15108 21480
rect 15160 21468 15166 21480
rect 15381 21471 15439 21477
rect 15381 21470 15393 21471
rect 15304 21468 15393 21470
rect 15160 21442 15393 21468
rect 15160 21440 15332 21442
rect 15160 21428 15166 21440
rect 15381 21437 15393 21442
rect 15427 21437 15439 21471
rect 15381 21431 15439 21437
rect 16761 21471 16819 21477
rect 16761 21437 16773 21471
rect 16807 21468 16819 21471
rect 16942 21468 16948 21480
rect 16807 21440 16948 21468
rect 16807 21437 16819 21440
rect 16761 21431 16819 21437
rect 16942 21428 16948 21440
rect 17000 21428 17006 21480
rect 18138 21428 18144 21480
rect 18196 21428 18202 21480
rect 19518 21428 19524 21480
rect 19576 21428 19582 21480
rect 19702 21477 19708 21480
rect 19675 21471 19708 21477
rect 19675 21437 19687 21471
rect 19760 21468 19766 21480
rect 20898 21468 20904 21480
rect 19760 21440 20904 21468
rect 19675 21431 19708 21437
rect 19702 21428 19708 21431
rect 19760 21428 19766 21440
rect 20898 21428 20904 21440
rect 20956 21428 20962 21480
rect 21358 21428 21364 21480
rect 21416 21428 21422 21480
rect 21468 21477 21496 21508
rect 21453 21471 21511 21477
rect 21453 21437 21465 21471
rect 21499 21437 21511 21471
rect 21453 21431 21511 21437
rect 21545 21471 21603 21477
rect 21545 21437 21557 21471
rect 21591 21468 21603 21471
rect 21634 21468 21640 21480
rect 21591 21440 21640 21468
rect 21591 21437 21603 21440
rect 21545 21431 21603 21437
rect 21634 21428 21640 21440
rect 21692 21428 21698 21480
rect 21821 21471 21879 21477
rect 21821 21437 21833 21471
rect 21867 21468 21879 21471
rect 21910 21468 21916 21480
rect 21867 21440 21916 21468
rect 21867 21437 21879 21440
rect 21821 21431 21879 21437
rect 21910 21428 21916 21440
rect 21968 21428 21974 21480
rect 15286 21400 15292 21412
rect 15028 21372 15292 21400
rect 15286 21360 15292 21372
rect 15344 21360 15350 21412
rect 16022 21360 16028 21412
rect 16080 21360 16086 21412
rect 16209 21403 16267 21409
rect 16209 21369 16221 21403
rect 16255 21369 16267 21403
rect 16209 21363 16267 21369
rect 13464 21304 14688 21332
rect 15105 21335 15163 21341
rect 15105 21301 15117 21335
rect 15151 21332 15163 21335
rect 15562 21332 15568 21344
rect 15151 21304 15568 21332
rect 15151 21301 15163 21304
rect 15105 21295 15163 21301
rect 15562 21292 15568 21304
rect 15620 21292 15626 21344
rect 15749 21335 15807 21341
rect 15749 21301 15761 21335
rect 15795 21332 15807 21335
rect 15930 21332 15936 21344
rect 15795 21304 15936 21332
rect 15795 21301 15807 21304
rect 15749 21295 15807 21301
rect 15930 21292 15936 21304
rect 15988 21332 15994 21344
rect 16224 21332 16252 21363
rect 17218 21360 17224 21412
rect 17276 21360 17282 21412
rect 17681 21403 17739 21409
rect 17681 21369 17693 21403
rect 17727 21369 17739 21403
rect 17681 21363 17739 21369
rect 15988 21304 16252 21332
rect 15988 21292 15994 21304
rect 17034 21292 17040 21344
rect 17092 21332 17098 21344
rect 17129 21335 17187 21341
rect 17129 21332 17141 21335
rect 17092 21304 17141 21332
rect 17092 21292 17098 21304
rect 17129 21301 17141 21304
rect 17175 21332 17187 21335
rect 17421 21335 17479 21341
rect 17421 21332 17433 21335
rect 17175 21304 17433 21332
rect 17175 21301 17187 21304
rect 17129 21295 17187 21301
rect 17421 21301 17433 21304
rect 17467 21301 17479 21335
rect 17421 21295 17479 21301
rect 17589 21335 17647 21341
rect 17589 21301 17601 21335
rect 17635 21332 17647 21335
rect 17696 21332 17724 21363
rect 17862 21360 17868 21412
rect 17920 21400 17926 21412
rect 18417 21403 18475 21409
rect 18417 21400 18429 21403
rect 17920 21372 18429 21400
rect 17920 21360 17926 21372
rect 18417 21369 18429 21372
rect 18463 21369 18475 21403
rect 18417 21363 18475 21369
rect 19242 21360 19248 21412
rect 19300 21400 19306 21412
rect 20441 21403 20499 21409
rect 19300 21372 20024 21400
rect 19300 21360 19306 21372
rect 17635 21304 17724 21332
rect 17635 21301 17647 21304
rect 17589 21295 17647 21301
rect 18046 21292 18052 21344
rect 18104 21292 18110 21344
rect 18230 21292 18236 21344
rect 18288 21292 18294 21344
rect 19426 21292 19432 21344
rect 19484 21332 19490 21344
rect 19889 21335 19947 21341
rect 19889 21332 19901 21335
rect 19484 21304 19901 21332
rect 19484 21292 19490 21304
rect 19889 21301 19901 21304
rect 19935 21301 19947 21335
rect 19996 21332 20024 21372
rect 20441 21369 20453 21403
rect 20487 21400 20499 21403
rect 20714 21400 20720 21412
rect 20487 21372 20720 21400
rect 20487 21369 20499 21372
rect 20441 21363 20499 21369
rect 20714 21360 20720 21372
rect 20772 21360 20778 21412
rect 20993 21403 21051 21409
rect 20993 21369 21005 21403
rect 21039 21400 21051 21403
rect 21726 21400 21732 21412
rect 21039 21372 21732 21400
rect 21039 21369 21051 21372
rect 20993 21363 21051 21369
rect 21726 21360 21732 21372
rect 21784 21360 21790 21412
rect 20898 21332 20904 21344
rect 19996 21304 20904 21332
rect 19889 21295 19947 21301
rect 20898 21292 20904 21304
rect 20956 21292 20962 21344
rect 21450 21292 21456 21344
rect 21508 21332 21514 21344
rect 21637 21335 21695 21341
rect 21637 21332 21649 21335
rect 21508 21304 21649 21332
rect 21508 21292 21514 21304
rect 21637 21301 21649 21304
rect 21683 21301 21695 21335
rect 21637 21295 21695 21301
rect 552 21242 23368 21264
rect 552 21190 4322 21242
rect 4374 21190 4386 21242
rect 4438 21190 4450 21242
rect 4502 21190 4514 21242
rect 4566 21190 4578 21242
rect 4630 21190 23368 21242
rect 552 21168 23368 21190
rect 7745 21131 7803 21137
rect 5276 21100 7604 21128
rect 4522 21020 4528 21072
rect 4580 21020 4586 21072
rect 5276 21060 5304 21100
rect 4908 21032 5304 21060
rect 4246 20952 4252 21004
rect 4304 20992 4310 21004
rect 4433 20995 4491 21001
rect 4433 20992 4445 20995
rect 4304 20964 4445 20992
rect 4304 20952 4310 20964
rect 4433 20961 4445 20964
rect 4479 20992 4491 20995
rect 4908 20992 4936 21032
rect 7098 21020 7104 21072
rect 7156 21060 7162 21072
rect 7576 21060 7604 21100
rect 7745 21097 7757 21131
rect 7791 21128 7803 21131
rect 9766 21128 9772 21140
rect 7791 21100 9772 21128
rect 7791 21097 7803 21100
rect 7745 21091 7803 21097
rect 9766 21088 9772 21100
rect 9824 21088 9830 21140
rect 9953 21131 10011 21137
rect 9953 21097 9965 21131
rect 9999 21128 10011 21131
rect 10686 21128 10692 21140
rect 9999 21100 10692 21128
rect 9999 21097 10011 21100
rect 9953 21091 10011 21097
rect 10686 21088 10692 21100
rect 10744 21088 10750 21140
rect 14182 21128 14188 21140
rect 10796 21100 14188 21128
rect 8297 21063 8355 21069
rect 8297 21060 8309 21063
rect 7156 21032 7512 21060
rect 7576 21032 8309 21060
rect 7156 21020 7162 21032
rect 4479 20964 4936 20992
rect 4985 20995 5043 21001
rect 4479 20961 4491 20964
rect 4433 20955 4491 20961
rect 4985 20961 4997 20995
rect 5031 20992 5043 20995
rect 5074 20992 5080 21004
rect 5031 20964 5080 20992
rect 5031 20961 5043 20964
rect 4985 20955 5043 20961
rect 5074 20952 5080 20964
rect 5132 20992 5138 21004
rect 5132 20964 6408 20992
rect 5132 20952 5138 20964
rect 6380 20936 6408 20964
rect 7190 20952 7196 21004
rect 7248 20952 7254 21004
rect 7285 20995 7343 21001
rect 7285 20961 7297 20995
rect 7331 20992 7343 20995
rect 7374 20992 7380 21004
rect 7331 20964 7380 20992
rect 7331 20961 7343 20964
rect 7285 20955 7343 20961
rect 7374 20952 7380 20964
rect 7432 20952 7438 21004
rect 7484 21001 7512 21032
rect 8297 21029 8309 21032
rect 8343 21060 8355 21063
rect 8662 21060 8668 21072
rect 8343 21032 8668 21060
rect 8343 21029 8355 21032
rect 8297 21023 8355 21029
rect 8662 21020 8668 21032
rect 8720 21020 8726 21072
rect 9033 21063 9091 21069
rect 9033 21029 9045 21063
rect 9079 21060 9091 21063
rect 9079 21032 9904 21060
rect 9079 21029 9091 21032
rect 9033 21023 9091 21029
rect 7469 20995 7527 21001
rect 7469 20961 7481 20995
rect 7515 20961 7527 20995
rect 7469 20955 7527 20961
rect 7558 20952 7564 21004
rect 7616 20952 7622 21004
rect 8202 20952 8208 21004
rect 8260 20952 8266 21004
rect 8478 20952 8484 21004
rect 8536 20992 8542 21004
rect 8938 20992 8944 21004
rect 8536 20964 8944 20992
rect 8536 20952 8542 20964
rect 8938 20952 8944 20964
rect 8996 20952 9002 21004
rect 9122 20952 9128 21004
rect 9180 20952 9186 21004
rect 9214 20952 9220 21004
rect 9272 20952 9278 21004
rect 9306 20952 9312 21004
rect 9364 20992 9370 21004
rect 9876 21001 9904 21032
rect 10134 21020 10140 21072
rect 10192 21060 10198 21072
rect 10796 21060 10824 21100
rect 14182 21088 14188 21100
rect 14240 21088 14246 21140
rect 15010 21128 15016 21140
rect 14752 21100 15016 21128
rect 14752 21060 14780 21100
rect 15010 21088 15016 21100
rect 15068 21088 15074 21140
rect 15562 21088 15568 21140
rect 15620 21128 15626 21140
rect 16853 21131 16911 21137
rect 16853 21128 16865 21131
rect 15620 21100 16865 21128
rect 15620 21088 15626 21100
rect 16853 21097 16865 21100
rect 16899 21128 16911 21131
rect 17218 21128 17224 21140
rect 16899 21100 17224 21128
rect 16899 21097 16911 21100
rect 16853 21091 16911 21097
rect 17218 21088 17224 21100
rect 17276 21088 17282 21140
rect 10192 21032 10824 21060
rect 12406 21032 14780 21060
rect 10192 21020 10198 21032
rect 9401 20995 9459 21001
rect 9401 20992 9413 20995
rect 9364 20964 9413 20992
rect 9364 20952 9370 20964
rect 9401 20961 9413 20964
rect 9447 20961 9459 20995
rect 9401 20955 9459 20961
rect 9861 20995 9919 21001
rect 9861 20961 9873 20995
rect 9907 20961 9919 20995
rect 9861 20955 9919 20961
rect 10042 20952 10048 21004
rect 10100 20952 10106 21004
rect 12250 20952 12256 21004
rect 12308 20952 12314 21004
rect 6362 20884 6368 20936
rect 6420 20924 6426 20936
rect 8220 20924 8248 20952
rect 6420 20896 8248 20924
rect 9137 20924 9165 20952
rect 12406 20924 12434 21032
rect 14826 21020 14832 21072
rect 14884 21060 14890 21072
rect 15473 21063 15531 21069
rect 14884 21032 14964 21060
rect 14884 21020 14890 21032
rect 12713 20995 12771 21001
rect 12713 20961 12725 20995
rect 12759 20992 12771 20995
rect 12802 20992 12808 21004
rect 12759 20964 12808 20992
rect 12759 20961 12771 20964
rect 12713 20955 12771 20961
rect 12802 20952 12808 20964
rect 12860 20952 12866 21004
rect 13078 20952 13084 21004
rect 13136 20952 13142 21004
rect 13265 20995 13323 21001
rect 13265 20961 13277 20995
rect 13311 20961 13323 20995
rect 13265 20955 13323 20961
rect 9137 20896 12434 20924
rect 12621 20927 12679 20933
rect 6420 20884 6426 20896
rect 12621 20893 12633 20927
rect 12667 20924 12679 20927
rect 13280 20924 13308 20955
rect 14734 20952 14740 21004
rect 14792 20952 14798 21004
rect 14936 21001 14964 21032
rect 15473 21029 15485 21063
rect 15519 21060 15531 21063
rect 16022 21060 16028 21072
rect 15519 21032 16028 21060
rect 15519 21029 15531 21032
rect 15473 21023 15531 21029
rect 14921 20995 14979 21001
rect 14921 20961 14933 20995
rect 14967 20961 14979 20995
rect 14921 20955 14979 20961
rect 15381 20995 15439 21001
rect 15381 20961 15393 20995
rect 15427 20961 15439 20995
rect 15381 20955 15439 20961
rect 12667 20896 13308 20924
rect 12667 20893 12679 20896
rect 12621 20887 12679 20893
rect 8665 20859 8723 20865
rect 8665 20825 8677 20859
rect 8711 20856 8723 20859
rect 10686 20856 10692 20868
rect 8711 20828 10692 20856
rect 8711 20825 8723 20828
rect 8665 20819 8723 20825
rect 10686 20816 10692 20828
rect 10744 20816 10750 20868
rect 13280 20856 13308 20896
rect 14093 20927 14151 20933
rect 14093 20893 14105 20927
rect 14139 20924 14151 20927
rect 14182 20924 14188 20936
rect 14139 20896 14188 20924
rect 14139 20893 14151 20896
rect 14093 20887 14151 20893
rect 14182 20884 14188 20896
rect 14240 20884 14246 20936
rect 14829 20927 14887 20933
rect 14829 20893 14841 20927
rect 14875 20924 14887 20927
rect 15396 20924 15424 20955
rect 15562 20952 15568 21004
rect 15620 20952 15626 21004
rect 15764 21001 15792 21032
rect 16022 21020 16028 21032
rect 16080 21020 16086 21072
rect 17034 21020 17040 21072
rect 17092 21020 17098 21072
rect 15749 20995 15807 21001
rect 15749 20961 15761 20995
rect 15795 20961 15807 20995
rect 15749 20955 15807 20961
rect 15930 20952 15936 21004
rect 15988 20952 15994 21004
rect 16393 20995 16451 21001
rect 16393 20961 16405 20995
rect 16439 20961 16451 20995
rect 16393 20955 16451 20961
rect 16577 20995 16635 21001
rect 16577 20961 16589 20995
rect 16623 20992 16635 20995
rect 16758 20992 16764 21004
rect 16623 20964 16764 20992
rect 16623 20961 16635 20964
rect 16577 20955 16635 20961
rect 14875 20896 15424 20924
rect 15841 20927 15899 20933
rect 14875 20893 14887 20896
rect 14829 20887 14887 20893
rect 15841 20893 15853 20927
rect 15887 20924 15899 20927
rect 16408 20924 16436 20955
rect 16758 20952 16764 20964
rect 16816 20952 16822 21004
rect 17405 20995 17463 21001
rect 17405 20961 17417 20995
rect 17451 20992 17463 20995
rect 18230 20992 18236 21004
rect 17451 20964 18236 20992
rect 17451 20961 17463 20964
rect 17405 20955 17463 20961
rect 17420 20924 17448 20955
rect 18230 20952 18236 20964
rect 18288 20952 18294 21004
rect 19518 20952 19524 21004
rect 19576 21001 19582 21004
rect 19576 20995 19609 21001
rect 19597 20961 19609 20995
rect 19576 20955 19609 20961
rect 19576 20952 19582 20955
rect 19702 20952 19708 21004
rect 19760 20952 19766 21004
rect 20622 20952 20628 21004
rect 20680 20992 20686 21004
rect 21637 20995 21695 21001
rect 21637 20992 21649 20995
rect 20680 20964 21649 20992
rect 20680 20952 20686 20964
rect 21637 20961 21649 20964
rect 21683 20961 21695 20995
rect 21637 20955 21695 20961
rect 21726 20952 21732 21004
rect 21784 20992 21790 21004
rect 22373 20995 22431 21001
rect 22373 20992 22385 20995
rect 21784 20964 22385 20992
rect 21784 20952 21790 20964
rect 22373 20961 22385 20964
rect 22419 20961 22431 20995
rect 22373 20955 22431 20961
rect 15887 20896 16436 20924
rect 16960 20896 17448 20924
rect 17497 20927 17555 20933
rect 15887 20893 15899 20896
rect 15841 20887 15899 20893
rect 16298 20856 16304 20868
rect 13280 20828 16304 20856
rect 16298 20816 16304 20828
rect 16356 20856 16362 20868
rect 16960 20856 16988 20896
rect 17497 20893 17509 20927
rect 17543 20924 17555 20927
rect 18046 20924 18052 20936
rect 17543 20896 18052 20924
rect 17543 20893 17555 20896
rect 17497 20887 17555 20893
rect 18046 20884 18052 20896
rect 18104 20884 18110 20936
rect 21453 20927 21511 20933
rect 21453 20893 21465 20927
rect 21499 20893 21511 20927
rect 21453 20887 21511 20893
rect 16356 20828 16988 20856
rect 17037 20859 17095 20865
rect 16356 20816 16362 20828
rect 17037 20825 17049 20859
rect 17083 20856 17095 20859
rect 17862 20856 17868 20868
rect 17083 20828 17868 20856
rect 17083 20825 17095 20828
rect 17037 20819 17095 20825
rect 17862 20816 17868 20828
rect 17920 20816 17926 20868
rect 20990 20816 20996 20868
rect 21048 20856 21054 20868
rect 21468 20856 21496 20887
rect 21542 20884 21548 20936
rect 21600 20884 21606 20936
rect 22094 20856 22100 20868
rect 21048 20828 21404 20856
rect 21468 20828 22100 20856
rect 21048 20816 21054 20828
rect 9030 20748 9036 20800
rect 9088 20788 9094 20800
rect 9309 20791 9367 20797
rect 9309 20788 9321 20791
rect 9088 20760 9321 20788
rect 9088 20748 9094 20760
rect 9309 20757 9321 20760
rect 9355 20757 9367 20791
rect 9309 20751 9367 20757
rect 9398 20748 9404 20800
rect 9456 20788 9462 20800
rect 11146 20788 11152 20800
rect 9456 20760 11152 20788
rect 9456 20748 9462 20760
rect 11146 20748 11152 20760
rect 11204 20748 11210 20800
rect 12802 20748 12808 20800
rect 12860 20788 12866 20800
rect 12897 20791 12955 20797
rect 12897 20788 12909 20791
rect 12860 20760 12909 20788
rect 12860 20748 12866 20760
rect 12897 20757 12909 20760
rect 12943 20757 12955 20791
rect 12897 20751 12955 20757
rect 16206 20748 16212 20800
rect 16264 20748 16270 20800
rect 17770 20748 17776 20800
rect 17828 20748 17834 20800
rect 19521 20791 19579 20797
rect 19521 20757 19533 20791
rect 19567 20788 19579 20791
rect 19610 20788 19616 20800
rect 19567 20760 19616 20788
rect 19567 20757 19579 20760
rect 19521 20751 19579 20757
rect 19610 20748 19616 20760
rect 19668 20748 19674 20800
rect 21266 20748 21272 20800
rect 21324 20748 21330 20800
rect 21376 20788 21404 20828
rect 22094 20816 22100 20828
rect 22152 20816 22158 20868
rect 21542 20788 21548 20800
rect 21376 20760 21548 20788
rect 21542 20748 21548 20760
rect 21600 20788 21606 20800
rect 21913 20791 21971 20797
rect 21913 20788 21925 20791
rect 21600 20760 21925 20788
rect 21600 20748 21606 20760
rect 21913 20757 21925 20760
rect 21959 20757 21971 20791
rect 21913 20751 21971 20757
rect 552 20698 23368 20720
rect 552 20646 3662 20698
rect 3714 20646 3726 20698
rect 3778 20646 3790 20698
rect 3842 20646 3854 20698
rect 3906 20646 3918 20698
rect 3970 20646 23368 20698
rect 552 20624 23368 20646
rect 4522 20544 4528 20596
rect 4580 20584 4586 20596
rect 5258 20584 5264 20596
rect 4580 20556 5264 20584
rect 4580 20544 4586 20556
rect 5258 20544 5264 20556
rect 5316 20544 5322 20596
rect 9217 20587 9275 20593
rect 9217 20553 9229 20587
rect 9263 20584 9275 20587
rect 10042 20584 10048 20596
rect 9263 20556 10048 20584
rect 9263 20553 9275 20556
rect 9217 20547 9275 20553
rect 10042 20544 10048 20556
rect 10100 20584 10106 20596
rect 10962 20584 10968 20596
rect 10100 20556 10968 20584
rect 10100 20544 10106 20556
rect 10962 20544 10968 20556
rect 11020 20544 11026 20596
rect 20809 20587 20867 20593
rect 20809 20553 20821 20587
rect 20855 20584 20867 20587
rect 21085 20587 21143 20593
rect 21085 20584 21097 20587
rect 20855 20556 21097 20584
rect 20855 20553 20867 20556
rect 20809 20547 20867 20553
rect 21085 20553 21097 20556
rect 21131 20553 21143 20587
rect 21085 20547 21143 20553
rect 21545 20587 21603 20593
rect 21545 20553 21557 20587
rect 21591 20553 21603 20587
rect 21545 20547 21603 20553
rect 4709 20519 4767 20525
rect 4709 20485 4721 20519
rect 4755 20516 4767 20519
rect 4798 20516 4804 20528
rect 4755 20488 4804 20516
rect 4755 20485 4767 20488
rect 4709 20479 4767 20485
rect 4798 20476 4804 20488
rect 4856 20476 4862 20528
rect 21450 20516 21456 20528
rect 20548 20488 21456 20516
rect 4433 20451 4491 20457
rect 4433 20417 4445 20451
rect 4479 20448 4491 20451
rect 6270 20448 6276 20460
rect 4479 20420 6276 20448
rect 4479 20417 4491 20420
rect 4433 20411 4491 20417
rect 4341 20383 4399 20389
rect 4341 20349 4353 20383
rect 4387 20380 4399 20383
rect 4614 20380 4620 20392
rect 4387 20352 4620 20380
rect 4387 20349 4399 20352
rect 4341 20343 4399 20349
rect 4614 20340 4620 20352
rect 4672 20340 4678 20392
rect 4801 20383 4859 20389
rect 4801 20349 4813 20383
rect 4847 20349 4859 20383
rect 4801 20343 4859 20349
rect 4062 20272 4068 20324
rect 4120 20312 4126 20324
rect 4816 20312 4844 20343
rect 4982 20340 4988 20392
rect 5040 20340 5046 20392
rect 5258 20340 5264 20392
rect 5316 20340 5322 20392
rect 5368 20389 5396 20420
rect 6270 20408 6276 20420
rect 6328 20408 6334 20460
rect 5353 20383 5411 20389
rect 5353 20349 5365 20383
rect 5399 20380 5411 20383
rect 5399 20352 5433 20380
rect 5399 20349 5411 20352
rect 5353 20343 5411 20349
rect 5534 20340 5540 20392
rect 5592 20380 5598 20392
rect 7374 20380 7380 20392
rect 5592 20352 7380 20380
rect 5592 20340 5598 20352
rect 7374 20340 7380 20352
rect 7432 20340 7438 20392
rect 9030 20340 9036 20392
rect 9088 20380 9094 20392
rect 9217 20383 9275 20389
rect 9217 20380 9229 20383
rect 9088 20352 9229 20380
rect 9088 20340 9094 20352
rect 9217 20349 9229 20352
rect 9263 20349 9275 20383
rect 9217 20343 9275 20349
rect 9401 20383 9459 20389
rect 9401 20349 9413 20383
rect 9447 20380 9459 20383
rect 9582 20380 9588 20392
rect 9447 20352 9588 20380
rect 9447 20349 9459 20352
rect 9401 20343 9459 20349
rect 9582 20340 9588 20352
rect 9640 20380 9646 20392
rect 15102 20380 15108 20392
rect 9640 20352 15108 20380
rect 9640 20340 9646 20352
rect 15102 20340 15108 20352
rect 15160 20380 15166 20392
rect 16666 20380 16672 20392
rect 15160 20352 16672 20380
rect 15160 20340 15166 20352
rect 16666 20340 16672 20352
rect 16724 20340 16730 20392
rect 19426 20340 19432 20392
rect 19484 20340 19490 20392
rect 19610 20340 19616 20392
rect 19668 20340 19674 20392
rect 20438 20340 20444 20392
rect 20496 20380 20502 20392
rect 20548 20389 20576 20488
rect 21450 20476 21456 20488
rect 21508 20516 21514 20528
rect 21560 20516 21588 20547
rect 21508 20488 21588 20516
rect 21508 20476 21514 20488
rect 20622 20408 20628 20460
rect 20680 20448 20686 20460
rect 20680 20420 21680 20448
rect 20680 20408 20686 20420
rect 20533 20383 20591 20389
rect 20533 20380 20545 20383
rect 20496 20352 20545 20380
rect 20496 20340 20502 20352
rect 20533 20349 20545 20352
rect 20579 20349 20591 20383
rect 20533 20343 20591 20349
rect 20714 20340 20720 20392
rect 20772 20380 20778 20392
rect 21085 20383 21143 20389
rect 21085 20380 21097 20383
rect 20772 20352 21097 20380
rect 20772 20340 20778 20352
rect 21085 20349 21097 20352
rect 21131 20349 21143 20383
rect 21085 20343 21143 20349
rect 21269 20383 21327 20389
rect 21269 20349 21281 20383
rect 21315 20349 21327 20383
rect 21269 20343 21327 20349
rect 4120 20284 4844 20312
rect 4120 20272 4126 20284
rect 4890 20272 4896 20324
rect 4948 20312 4954 20324
rect 14734 20312 14740 20324
rect 4948 20284 14740 20312
rect 4948 20272 4954 20284
rect 14734 20272 14740 20284
rect 14792 20272 14798 20324
rect 19444 20312 19472 20340
rect 20622 20312 20628 20324
rect 19444 20284 20628 20312
rect 20622 20272 20628 20284
rect 20680 20272 20686 20324
rect 20809 20315 20867 20321
rect 20809 20281 20821 20315
rect 20855 20312 20867 20315
rect 20990 20312 20996 20324
rect 20855 20284 20996 20312
rect 20855 20281 20867 20284
rect 20809 20275 20867 20281
rect 20990 20272 20996 20284
rect 21048 20272 21054 20324
rect 5721 20247 5779 20253
rect 5721 20213 5733 20247
rect 5767 20244 5779 20247
rect 6730 20244 6736 20256
rect 5767 20216 6736 20244
rect 5767 20213 5779 20216
rect 5721 20207 5779 20213
rect 6730 20204 6736 20216
rect 6788 20204 6794 20256
rect 19150 20204 19156 20256
rect 19208 20244 19214 20256
rect 19429 20247 19487 20253
rect 19429 20244 19441 20247
rect 19208 20216 19441 20244
rect 19208 20204 19214 20216
rect 19429 20213 19441 20216
rect 19475 20213 19487 20247
rect 19429 20207 19487 20213
rect 20714 20204 20720 20256
rect 20772 20244 20778 20256
rect 20901 20247 20959 20253
rect 20901 20244 20913 20247
rect 20772 20216 20913 20244
rect 20772 20204 20778 20216
rect 20901 20213 20913 20216
rect 20947 20213 20959 20247
rect 21284 20244 21312 20343
rect 21542 20321 21548 20324
rect 21529 20315 21548 20321
rect 21529 20281 21541 20315
rect 21529 20275 21548 20281
rect 21542 20272 21548 20275
rect 21600 20272 21606 20324
rect 21652 20312 21680 20420
rect 21729 20315 21787 20321
rect 21729 20312 21741 20315
rect 21652 20284 21741 20312
rect 21729 20281 21741 20284
rect 21775 20281 21787 20315
rect 21729 20275 21787 20281
rect 21361 20247 21419 20253
rect 21361 20244 21373 20247
rect 21284 20216 21373 20244
rect 20901 20207 20959 20213
rect 21361 20213 21373 20216
rect 21407 20213 21419 20247
rect 21361 20207 21419 20213
rect 552 20154 23368 20176
rect 552 20102 4322 20154
rect 4374 20102 4386 20154
rect 4438 20102 4450 20154
rect 4502 20102 4514 20154
rect 4566 20102 4578 20154
rect 4630 20102 23368 20154
rect 552 20080 23368 20102
rect 5074 20040 5080 20052
rect 4356 20012 5080 20040
rect 2866 19932 2872 19984
rect 2924 19972 2930 19984
rect 2924 19944 3004 19972
rect 2924 19932 2930 19944
rect 2774 19864 2780 19916
rect 2832 19864 2838 19916
rect 2976 19913 3004 19944
rect 3326 19932 3332 19984
rect 3384 19972 3390 19984
rect 4062 19972 4068 19984
rect 3384 19944 4068 19972
rect 3384 19932 3390 19944
rect 4062 19932 4068 19944
rect 4120 19972 4126 19984
rect 4356 19981 4384 20012
rect 5074 20000 5080 20012
rect 5132 20000 5138 20052
rect 21266 20000 21272 20052
rect 21324 20000 21330 20052
rect 4157 19975 4215 19981
rect 4157 19972 4169 19975
rect 4120 19944 4169 19972
rect 4120 19932 4126 19944
rect 4157 19941 4169 19944
rect 4203 19941 4215 19975
rect 4157 19935 4215 19941
rect 4341 19975 4399 19981
rect 4341 19941 4353 19975
rect 4387 19941 4399 19975
rect 4341 19935 4399 19941
rect 4801 19975 4859 19981
rect 4801 19941 4813 19975
rect 4847 19972 4859 19975
rect 4982 19972 4988 19984
rect 4847 19944 4988 19972
rect 4847 19941 4859 19944
rect 4801 19935 4859 19941
rect 4982 19932 4988 19944
rect 5040 19972 5046 19984
rect 5353 19975 5411 19981
rect 5353 19972 5365 19975
rect 5040 19944 5365 19972
rect 5040 19932 5046 19944
rect 5353 19941 5365 19944
rect 5399 19941 5411 19975
rect 5353 19935 5411 19941
rect 2961 19907 3019 19913
rect 2961 19873 2973 19907
rect 3007 19873 3019 19907
rect 2961 19867 3019 19873
rect 3418 19864 3424 19916
rect 3476 19904 3482 19916
rect 3513 19907 3571 19913
rect 3513 19904 3525 19907
rect 3476 19876 3525 19904
rect 3476 19864 3482 19876
rect 3513 19873 3525 19876
rect 3559 19873 3571 19907
rect 3513 19867 3571 19873
rect 4525 19907 4583 19913
rect 4525 19873 4537 19907
rect 4571 19904 4583 19907
rect 4709 19907 4767 19913
rect 4709 19904 4721 19907
rect 4571 19876 4721 19904
rect 4571 19873 4583 19876
rect 4525 19867 4583 19873
rect 4709 19873 4721 19876
rect 4755 19873 4767 19907
rect 4709 19867 4767 19873
rect 4890 19864 4896 19916
rect 4948 19864 4954 19916
rect 5169 19907 5227 19913
rect 5169 19873 5181 19907
rect 5215 19873 5227 19907
rect 5169 19867 5227 19873
rect 8481 19907 8539 19913
rect 8481 19873 8493 19907
rect 8527 19904 8539 19907
rect 8754 19904 8760 19916
rect 8527 19876 8760 19904
rect 8527 19873 8539 19876
rect 8481 19867 8539 19873
rect 2869 19839 2927 19845
rect 2869 19805 2881 19839
rect 2915 19805 2927 19839
rect 5184 19836 5212 19867
rect 8754 19864 8760 19876
rect 8812 19864 8818 19916
rect 9122 19864 9128 19916
rect 9180 19864 9186 19916
rect 9858 19864 9864 19916
rect 9916 19864 9922 19916
rect 11149 19907 11207 19913
rect 11149 19904 11161 19907
rect 10244 19876 11161 19904
rect 2869 19799 2927 19805
rect 4908 19808 5212 19836
rect 2884 19768 2912 19799
rect 4908 19780 4936 19808
rect 9490 19796 9496 19848
rect 9548 19836 9554 19848
rect 9769 19839 9827 19845
rect 9769 19836 9781 19839
rect 9548 19808 9781 19836
rect 9548 19796 9554 19808
rect 9769 19805 9781 19808
rect 9815 19805 9827 19839
rect 9769 19799 9827 19805
rect 2884 19740 3280 19768
rect 3252 19712 3280 19740
rect 4890 19728 4896 19780
rect 4948 19728 4954 19780
rect 10244 19777 10272 19876
rect 11149 19873 11161 19876
rect 11195 19904 11207 19907
rect 11238 19904 11244 19916
rect 11195 19876 11244 19904
rect 11195 19873 11207 19876
rect 11149 19867 11207 19873
rect 11238 19864 11244 19876
rect 11296 19864 11302 19916
rect 18690 19864 18696 19916
rect 18748 19904 18754 19916
rect 18877 19907 18935 19913
rect 18877 19904 18889 19907
rect 18748 19876 18889 19904
rect 18748 19864 18754 19876
rect 18877 19873 18889 19876
rect 18923 19873 18935 19907
rect 18877 19867 18935 19873
rect 19058 19864 19064 19916
rect 19116 19864 19122 19916
rect 19150 19864 19156 19916
rect 19208 19864 19214 19916
rect 19334 19864 19340 19916
rect 19392 19904 19398 19916
rect 20533 19907 20591 19913
rect 20533 19904 20545 19907
rect 19392 19876 20545 19904
rect 19392 19864 19398 19876
rect 20533 19873 20545 19876
rect 20579 19904 20591 19907
rect 20625 19907 20683 19913
rect 20625 19904 20637 19907
rect 20579 19876 20637 19904
rect 20579 19873 20591 19876
rect 20533 19867 20591 19873
rect 20625 19873 20637 19876
rect 20671 19873 20683 19907
rect 20625 19867 20683 19873
rect 20990 19864 20996 19916
rect 21048 19864 21054 19916
rect 21634 19864 21640 19916
rect 21692 19864 21698 19916
rect 11054 19796 11060 19848
rect 11112 19796 11118 19848
rect 21358 19796 21364 19848
rect 21416 19836 21422 19848
rect 21729 19839 21787 19845
rect 21729 19836 21741 19839
rect 21416 19808 21741 19836
rect 21416 19796 21422 19808
rect 21729 19805 21741 19808
rect 21775 19805 21787 19839
rect 21729 19799 21787 19805
rect 10229 19771 10287 19777
rect 10229 19737 10241 19771
rect 10275 19737 10287 19771
rect 10229 19731 10287 19737
rect 3142 19660 3148 19712
rect 3200 19660 3206 19712
rect 3234 19660 3240 19712
rect 3292 19700 3298 19712
rect 3329 19703 3387 19709
rect 3329 19700 3341 19703
rect 3292 19672 3341 19700
rect 3292 19660 3298 19672
rect 3329 19669 3341 19672
rect 3375 19669 3387 19703
rect 3329 19663 3387 19669
rect 5537 19703 5595 19709
rect 5537 19669 5549 19703
rect 5583 19700 5595 19703
rect 5994 19700 6000 19712
rect 5583 19672 6000 19700
rect 5583 19669 5595 19672
rect 5537 19663 5595 19669
rect 5994 19660 6000 19672
rect 6052 19660 6058 19712
rect 7650 19660 7656 19712
rect 7708 19660 7714 19712
rect 11514 19660 11520 19712
rect 11572 19660 11578 19712
rect 19153 19703 19211 19709
rect 19153 19669 19165 19703
rect 19199 19700 19211 19703
rect 19426 19700 19432 19712
rect 19199 19672 19432 19700
rect 19199 19669 19211 19672
rect 19153 19663 19211 19669
rect 19426 19660 19432 19672
rect 19484 19660 19490 19712
rect 19610 19660 19616 19712
rect 19668 19700 19674 19712
rect 20346 19700 20352 19712
rect 19668 19672 20352 19700
rect 19668 19660 19674 19672
rect 20346 19660 20352 19672
rect 20404 19660 20410 19712
rect 20530 19660 20536 19712
rect 20588 19700 20594 19712
rect 21913 19703 21971 19709
rect 21913 19700 21925 19703
rect 20588 19672 21925 19700
rect 20588 19660 20594 19672
rect 21913 19669 21925 19672
rect 21959 19669 21971 19703
rect 21913 19663 21971 19669
rect 552 19610 23368 19632
rect 552 19558 3662 19610
rect 3714 19558 3726 19610
rect 3778 19558 3790 19610
rect 3842 19558 3854 19610
rect 3906 19558 3918 19610
rect 3970 19558 23368 19610
rect 552 19536 23368 19558
rect 3881 19499 3939 19505
rect 3881 19465 3893 19499
rect 3927 19465 3939 19499
rect 3881 19459 3939 19465
rect 5261 19499 5319 19505
rect 5261 19465 5273 19499
rect 5307 19496 5319 19499
rect 5442 19496 5448 19508
rect 5307 19468 5448 19496
rect 5307 19465 5319 19468
rect 5261 19459 5319 19465
rect 2866 19388 2872 19440
rect 2924 19388 2930 19440
rect 3142 19388 3148 19440
rect 3200 19428 3206 19440
rect 3513 19431 3571 19437
rect 3513 19428 3525 19431
rect 3200 19400 3525 19428
rect 3200 19388 3206 19400
rect 3513 19397 3525 19400
rect 3559 19428 3571 19431
rect 3694 19428 3700 19440
rect 3559 19400 3700 19428
rect 3559 19397 3571 19400
rect 3513 19391 3571 19397
rect 3694 19388 3700 19400
rect 3752 19428 3758 19440
rect 3896 19428 3924 19459
rect 5442 19456 5448 19468
rect 5500 19496 5506 19508
rect 5813 19499 5871 19505
rect 5813 19496 5825 19499
rect 5500 19468 5825 19496
rect 5500 19456 5506 19468
rect 5813 19465 5825 19468
rect 5859 19465 5871 19499
rect 5813 19459 5871 19465
rect 6181 19499 6239 19505
rect 6181 19465 6193 19499
rect 6227 19496 6239 19499
rect 17037 19499 17095 19505
rect 6227 19468 15976 19496
rect 6227 19465 6239 19468
rect 6181 19459 6239 19465
rect 7190 19428 7196 19440
rect 3752 19400 3924 19428
rect 5736 19400 7196 19428
rect 3752 19388 3758 19400
rect 3053 19363 3111 19369
rect 3053 19329 3065 19363
rect 3099 19360 3111 19363
rect 3421 19363 3479 19369
rect 3421 19360 3433 19363
rect 3099 19332 3433 19360
rect 3099 19329 3111 19332
rect 3053 19323 3111 19329
rect 3421 19329 3433 19332
rect 3467 19329 3479 19363
rect 3973 19363 4031 19369
rect 3973 19360 3985 19363
rect 3421 19323 3479 19329
rect 3620 19332 3985 19360
rect 2593 19295 2651 19301
rect 2593 19261 2605 19295
rect 2639 19292 2651 19295
rect 2774 19292 2780 19304
rect 2639 19264 2780 19292
rect 2639 19261 2651 19264
rect 2593 19255 2651 19261
rect 2774 19252 2780 19264
rect 2832 19252 2838 19304
rect 3326 19252 3332 19304
rect 3384 19252 3390 19304
rect 3436 19224 3464 19323
rect 3620 19304 3648 19332
rect 3973 19329 3985 19332
rect 4019 19329 4031 19363
rect 3973 19323 4031 19329
rect 4890 19320 4896 19372
rect 4948 19320 4954 19372
rect 5736 19369 5764 19400
rect 7190 19388 7196 19400
rect 7248 19428 7254 19440
rect 7650 19428 7656 19440
rect 7248 19400 7656 19428
rect 7248 19388 7254 19400
rect 7650 19388 7656 19400
rect 7708 19388 7714 19440
rect 12345 19431 12403 19437
rect 12345 19397 12357 19431
rect 12391 19397 12403 19431
rect 12345 19391 12403 19397
rect 5721 19363 5779 19369
rect 5721 19329 5733 19363
rect 5767 19329 5779 19363
rect 5721 19323 5779 19329
rect 6730 19320 6736 19372
rect 6788 19320 6794 19372
rect 7285 19363 7343 19369
rect 7285 19360 7297 19363
rect 7116 19332 7297 19360
rect 3602 19252 3608 19304
rect 3660 19252 3666 19304
rect 3881 19295 3939 19301
rect 3881 19261 3893 19295
rect 3927 19261 3939 19295
rect 3881 19255 3939 19261
rect 3510 19224 3516 19236
rect 3436 19196 3516 19224
rect 3510 19184 3516 19196
rect 3568 19224 3574 19236
rect 3896 19224 3924 19255
rect 4982 19252 4988 19304
rect 5040 19252 5046 19304
rect 5276 19264 5948 19292
rect 5276 19224 5304 19264
rect 3568 19196 3924 19224
rect 4172 19196 5304 19224
rect 5920 19224 5948 19264
rect 5994 19252 6000 19304
rect 6052 19252 6058 19304
rect 6641 19295 6699 19301
rect 6641 19261 6653 19295
rect 6687 19292 6699 19295
rect 7116 19292 7144 19332
rect 7285 19329 7297 19332
rect 7331 19360 7343 19363
rect 7374 19360 7380 19372
rect 7331 19332 7380 19360
rect 7331 19329 7343 19332
rect 7285 19323 7343 19329
rect 7374 19320 7380 19332
rect 7432 19320 7438 19372
rect 11514 19320 11520 19372
rect 11572 19360 11578 19372
rect 11885 19363 11943 19369
rect 11885 19360 11897 19363
rect 11572 19332 11897 19360
rect 11572 19320 11578 19332
rect 11885 19329 11897 19332
rect 11931 19360 11943 19363
rect 12158 19360 12164 19372
rect 11931 19332 12164 19360
rect 11931 19329 11943 19332
rect 11885 19323 11943 19329
rect 12158 19320 12164 19332
rect 12216 19320 12222 19372
rect 12360 19360 12388 19391
rect 13081 19363 13139 19369
rect 12360 19332 13032 19360
rect 13004 19304 13032 19332
rect 13081 19329 13093 19363
rect 13127 19329 13139 19363
rect 13081 19323 13139 19329
rect 6687 19264 7144 19292
rect 7193 19295 7251 19301
rect 6687 19261 6699 19264
rect 6641 19255 6699 19261
rect 7193 19261 7205 19295
rect 7239 19292 7251 19295
rect 8386 19292 8392 19304
rect 7239 19264 8392 19292
rect 7239 19261 7251 19264
rect 7193 19255 7251 19261
rect 8386 19252 8392 19264
rect 8444 19252 8450 19304
rect 8754 19252 8760 19304
rect 8812 19292 8818 19304
rect 10229 19295 10287 19301
rect 8812 19264 9674 19292
rect 8812 19252 8818 19264
rect 6917 19227 6975 19233
rect 5920 19196 6868 19224
rect 3568 19184 3574 19196
rect 3789 19159 3847 19165
rect 3789 19125 3801 19159
rect 3835 19156 3847 19159
rect 4172 19156 4200 19196
rect 3835 19128 4200 19156
rect 3835 19125 3847 19128
rect 3789 19119 3847 19125
rect 4246 19116 4252 19168
rect 4304 19116 4310 19168
rect 6270 19116 6276 19168
rect 6328 19116 6334 19168
rect 6840 19156 6868 19196
rect 6917 19193 6929 19227
rect 6963 19224 6975 19227
rect 9490 19224 9496 19236
rect 6963 19196 9496 19224
rect 6963 19193 6975 19196
rect 6917 19187 6975 19193
rect 9490 19184 9496 19196
rect 9548 19184 9554 19236
rect 9646 19224 9674 19264
rect 10229 19261 10241 19295
rect 10275 19292 10287 19295
rect 10275 19264 10548 19292
rect 10275 19261 10287 19264
rect 10229 19255 10287 19261
rect 9766 19224 9772 19236
rect 9646 19196 9772 19224
rect 9766 19184 9772 19196
rect 9824 19224 9830 19236
rect 10520 19224 10548 19264
rect 10686 19252 10692 19304
rect 10744 19252 10750 19304
rect 10962 19252 10968 19304
rect 11020 19292 11026 19304
rect 11977 19295 12035 19301
rect 11977 19292 11989 19295
rect 11020 19264 11989 19292
rect 11020 19252 11026 19264
rect 11977 19261 11989 19264
rect 12023 19261 12035 19295
rect 11977 19255 12035 19261
rect 12986 19252 12992 19304
rect 13044 19252 13050 19304
rect 13096 19292 13124 19323
rect 13170 19320 13176 19372
rect 13228 19360 13234 19372
rect 15948 19369 15976 19468
rect 17037 19465 17049 19499
rect 17083 19496 17095 19499
rect 17497 19499 17555 19505
rect 17497 19496 17509 19499
rect 17083 19468 17509 19496
rect 17083 19465 17095 19468
rect 17037 19459 17095 19465
rect 17497 19465 17509 19468
rect 17543 19496 17555 19499
rect 17586 19496 17592 19508
rect 17543 19468 17592 19496
rect 17543 19465 17555 19468
rect 17497 19459 17555 19465
rect 17586 19456 17592 19468
rect 17644 19456 17650 19508
rect 17604 19428 17632 19456
rect 17604 19400 18276 19428
rect 13357 19363 13415 19369
rect 13357 19360 13369 19363
rect 13228 19332 13369 19360
rect 13228 19320 13234 19332
rect 13357 19329 13369 19332
rect 13403 19329 13415 19363
rect 13357 19323 13415 19329
rect 15933 19363 15991 19369
rect 15933 19329 15945 19363
rect 15979 19360 15991 19363
rect 15979 19332 16528 19360
rect 15979 19329 15991 19332
rect 15933 19323 15991 19329
rect 13262 19292 13268 19304
rect 13096 19264 13268 19292
rect 13262 19252 13268 19264
rect 13320 19252 13326 19304
rect 16025 19295 16083 19301
rect 16025 19261 16037 19295
rect 16071 19292 16083 19295
rect 16206 19292 16212 19304
rect 16071 19264 16212 19292
rect 16071 19261 16083 19264
rect 16025 19255 16083 19261
rect 16206 19252 16212 19264
rect 16264 19252 16270 19304
rect 16500 19301 16528 19332
rect 17770 19320 17776 19372
rect 17828 19360 17834 19372
rect 18141 19363 18199 19369
rect 18141 19360 18153 19363
rect 17828 19332 18153 19360
rect 17828 19320 17834 19332
rect 18141 19329 18153 19332
rect 18187 19329 18199 19363
rect 18141 19323 18199 19329
rect 16485 19295 16543 19301
rect 16485 19261 16497 19295
rect 16531 19261 16543 19295
rect 16485 19255 16543 19261
rect 16578 19295 16636 19301
rect 16578 19261 16590 19295
rect 16624 19261 16636 19295
rect 16945 19295 17003 19301
rect 16945 19292 16957 19295
rect 16578 19255 16636 19261
rect 16684 19264 16957 19292
rect 10594 19224 10600 19236
rect 9824 19196 9890 19224
rect 10520 19196 10600 19224
rect 9824 19184 9830 19196
rect 10594 19184 10600 19196
rect 10652 19224 10658 19236
rect 15194 19224 15200 19236
rect 10652 19196 15200 19224
rect 10652 19184 10658 19196
rect 15194 19184 15200 19196
rect 15252 19184 15258 19236
rect 16224 19224 16252 19252
rect 16592 19224 16620 19255
rect 16224 19196 16620 19224
rect 7098 19156 7104 19168
rect 6840 19128 7104 19156
rect 7098 19116 7104 19128
rect 7156 19116 7162 19168
rect 7558 19116 7564 19168
rect 7616 19116 7622 19168
rect 16390 19116 16396 19168
rect 16448 19156 16454 19168
rect 16684 19156 16712 19264
rect 16945 19261 16957 19264
rect 16991 19261 17003 19295
rect 16945 19255 17003 19261
rect 17126 19252 17132 19304
rect 17184 19252 17190 19304
rect 17865 19295 17923 19301
rect 17865 19261 17877 19295
rect 17911 19261 17923 19295
rect 17865 19255 17923 19261
rect 16853 19227 16911 19233
rect 16853 19193 16865 19227
rect 16899 19224 16911 19227
rect 17310 19224 17316 19236
rect 16899 19196 17316 19224
rect 16899 19193 16911 19196
rect 16853 19187 16911 19193
rect 17310 19184 17316 19196
rect 17368 19184 17374 19236
rect 17529 19227 17587 19233
rect 17529 19193 17541 19227
rect 17575 19224 17587 19227
rect 17770 19224 17776 19236
rect 17575 19196 17776 19224
rect 17575 19193 17587 19196
rect 17529 19187 17587 19193
rect 17770 19184 17776 19196
rect 17828 19184 17834 19236
rect 17880 19224 17908 19255
rect 17954 19252 17960 19304
rect 18012 19252 18018 19304
rect 18049 19295 18107 19301
rect 18049 19261 18061 19295
rect 18095 19292 18107 19295
rect 18248 19292 18276 19400
rect 20346 19388 20352 19440
rect 20404 19428 20410 19440
rect 20404 19400 20944 19428
rect 20404 19388 20410 19400
rect 18325 19363 18383 19369
rect 18325 19329 18337 19363
rect 18371 19360 18383 19363
rect 18371 19332 18736 19360
rect 18371 19329 18383 19332
rect 18325 19323 18383 19329
rect 18708 19304 18736 19332
rect 19426 19320 19432 19372
rect 19484 19320 19490 19372
rect 18095 19264 18276 19292
rect 18095 19261 18107 19264
rect 18049 19255 18107 19261
rect 18690 19252 18696 19304
rect 18748 19252 18754 19304
rect 18969 19295 19027 19301
rect 18969 19261 18981 19295
rect 19015 19292 19027 19295
rect 19150 19292 19156 19304
rect 19015 19264 19156 19292
rect 19015 19261 19027 19264
rect 18969 19255 19027 19261
rect 19150 19252 19156 19264
rect 19208 19252 19214 19304
rect 19521 19295 19579 19301
rect 19521 19261 19533 19295
rect 19567 19261 19579 19295
rect 19521 19255 19579 19261
rect 18414 19224 18420 19236
rect 17880 19196 18420 19224
rect 18414 19184 18420 19196
rect 18472 19184 18478 19236
rect 19536 19224 19564 19255
rect 19610 19252 19616 19304
rect 19668 19252 19674 19304
rect 19702 19252 19708 19304
rect 19760 19252 19766 19304
rect 20346 19252 20352 19304
rect 20404 19252 20410 19304
rect 20530 19252 20536 19304
rect 20588 19252 20594 19304
rect 20717 19295 20775 19301
rect 20717 19261 20729 19295
rect 20763 19292 20775 19295
rect 20806 19292 20812 19304
rect 20763 19264 20812 19292
rect 20763 19261 20775 19264
rect 20717 19255 20775 19261
rect 20806 19252 20812 19264
rect 20864 19252 20870 19304
rect 20916 19292 20944 19400
rect 20993 19295 21051 19301
rect 20993 19292 21005 19295
rect 20916 19264 21005 19292
rect 20993 19261 21005 19264
rect 21039 19261 21051 19295
rect 20993 19255 21051 19261
rect 21082 19252 21088 19304
rect 21140 19252 21146 19304
rect 21358 19252 21364 19304
rect 21416 19252 21422 19304
rect 21450 19252 21456 19304
rect 21508 19252 21514 19304
rect 22278 19252 22284 19304
rect 22336 19252 22342 19304
rect 22370 19252 22376 19304
rect 22428 19252 22434 19304
rect 22554 19252 22560 19304
rect 22612 19252 22618 19304
rect 23014 19252 23020 19304
rect 23072 19252 23078 19304
rect 20438 19224 20444 19236
rect 19168 19196 20444 19224
rect 16448 19128 16712 19156
rect 17681 19159 17739 19165
rect 16448 19116 16454 19128
rect 17681 19125 17693 19159
rect 17727 19156 17739 19159
rect 18046 19156 18052 19168
rect 17727 19128 18052 19156
rect 17727 19125 17739 19128
rect 17681 19119 17739 19125
rect 18046 19116 18052 19128
rect 18104 19116 18110 19168
rect 18138 19116 18144 19168
rect 18196 19156 18202 19168
rect 18785 19159 18843 19165
rect 18785 19156 18797 19159
rect 18196 19128 18797 19156
rect 18196 19116 18202 19128
rect 18785 19125 18797 19128
rect 18831 19156 18843 19159
rect 19058 19156 19064 19168
rect 18831 19128 19064 19156
rect 18831 19125 18843 19128
rect 18785 19119 18843 19125
rect 19058 19116 19064 19128
rect 19116 19116 19122 19168
rect 19168 19165 19196 19196
rect 20438 19184 20444 19196
rect 20496 19184 20502 19236
rect 20625 19227 20683 19233
rect 20625 19193 20637 19227
rect 20671 19224 20683 19227
rect 21174 19224 21180 19236
rect 20671 19196 21180 19224
rect 20671 19193 20683 19196
rect 20625 19187 20683 19193
rect 21174 19184 21180 19196
rect 21232 19184 21238 19236
rect 21376 19224 21404 19252
rect 21376 19196 21496 19224
rect 19153 19159 19211 19165
rect 19153 19125 19165 19159
rect 19199 19125 19211 19159
rect 19153 19119 19211 19125
rect 19242 19116 19248 19168
rect 19300 19116 19306 19168
rect 20901 19159 20959 19165
rect 20901 19125 20913 19159
rect 20947 19156 20959 19159
rect 21358 19156 21364 19168
rect 20947 19128 21364 19156
rect 20947 19125 20959 19128
rect 20901 19119 20959 19125
rect 21358 19116 21364 19128
rect 21416 19116 21422 19168
rect 21468 19165 21496 19196
rect 21453 19159 21511 19165
rect 21453 19125 21465 19159
rect 21499 19125 21511 19159
rect 21453 19119 21511 19125
rect 21634 19116 21640 19168
rect 21692 19116 21698 19168
rect 552 19066 23368 19088
rect 552 19014 4322 19066
rect 4374 19014 4386 19066
rect 4438 19014 4450 19066
rect 4502 19014 4514 19066
rect 4566 19014 4578 19066
rect 4630 19014 23368 19066
rect 552 18992 23368 19014
rect 3237 18955 3295 18961
rect 3237 18921 3249 18955
rect 3283 18952 3295 18955
rect 3602 18952 3608 18964
rect 3283 18924 3608 18952
rect 3283 18921 3295 18924
rect 3237 18915 3295 18921
rect 3602 18912 3608 18924
rect 3660 18912 3666 18964
rect 4249 18955 4307 18961
rect 4249 18921 4261 18955
rect 4295 18952 4307 18955
rect 5258 18952 5264 18964
rect 4295 18924 5264 18952
rect 4295 18921 4307 18924
rect 4249 18915 4307 18921
rect 5258 18912 5264 18924
rect 5316 18912 5322 18964
rect 6365 18955 6423 18961
rect 6365 18921 6377 18955
rect 6411 18952 6423 18955
rect 6411 18924 12112 18952
rect 6411 18921 6423 18924
rect 6365 18915 6423 18921
rect 2774 18844 2780 18896
rect 2832 18844 2838 18896
rect 4433 18887 4491 18893
rect 4433 18884 4445 18887
rect 3620 18856 4445 18884
rect 3620 18825 3648 18856
rect 4433 18853 4445 18856
rect 4479 18884 4491 18887
rect 5534 18884 5540 18896
rect 4479 18856 5540 18884
rect 4479 18853 4491 18856
rect 4433 18847 4491 18853
rect 5534 18844 5540 18856
rect 5592 18844 5598 18896
rect 5629 18887 5687 18893
rect 5629 18853 5641 18887
rect 5675 18884 5687 18887
rect 5675 18856 6224 18884
rect 5675 18853 5687 18856
rect 5629 18847 5687 18853
rect 3605 18819 3663 18825
rect 3605 18785 3617 18819
rect 3651 18785 3663 18819
rect 3605 18779 3663 18785
rect 3694 18776 3700 18828
rect 3752 18776 3758 18828
rect 4154 18776 4160 18828
rect 4212 18776 4218 18828
rect 4982 18776 4988 18828
rect 5040 18776 5046 18828
rect 5997 18819 6055 18825
rect 5997 18785 6009 18819
rect 6043 18785 6055 18819
rect 6196 18816 6224 18856
rect 6270 18844 6276 18896
rect 6328 18884 6334 18896
rect 6733 18887 6791 18893
rect 6733 18884 6745 18887
rect 6328 18856 6745 18884
rect 6328 18844 6334 18856
rect 6733 18853 6745 18856
rect 6779 18853 6791 18887
rect 8021 18887 8079 18893
rect 6733 18847 6791 18853
rect 6840 18856 7972 18884
rect 6457 18819 6515 18825
rect 6457 18816 6469 18819
rect 6196 18788 6469 18816
rect 5997 18779 6055 18785
rect 6457 18785 6469 18788
rect 6503 18785 6515 18819
rect 6457 18779 6515 18785
rect 5074 18708 5080 18760
rect 5132 18708 5138 18760
rect 5442 18708 5448 18760
rect 5500 18748 5506 18760
rect 5905 18751 5963 18757
rect 5905 18748 5917 18751
rect 5500 18720 5917 18748
rect 5500 18708 5506 18720
rect 5905 18717 5917 18720
rect 5951 18717 5963 18751
rect 6012 18748 6040 18779
rect 6472 18748 6500 18779
rect 6638 18776 6644 18828
rect 6696 18776 6702 18828
rect 6840 18825 6868 18856
rect 6825 18819 6883 18825
rect 6825 18785 6837 18819
rect 6871 18785 6883 18819
rect 6825 18779 6883 18785
rect 7282 18776 7288 18828
rect 7340 18816 7346 18828
rect 7469 18819 7527 18825
rect 7469 18816 7481 18819
rect 7340 18788 7481 18816
rect 7340 18776 7346 18788
rect 7469 18785 7481 18788
rect 7515 18785 7527 18819
rect 7469 18779 7527 18785
rect 7837 18819 7895 18825
rect 7837 18785 7849 18819
rect 7883 18785 7895 18819
rect 7944 18816 7972 18856
rect 8021 18853 8033 18887
rect 8067 18884 8079 18887
rect 9030 18884 9036 18896
rect 8067 18856 9036 18884
rect 8067 18853 8079 18856
rect 8021 18847 8079 18853
rect 9030 18844 9036 18856
rect 9088 18844 9094 18896
rect 10686 18884 10692 18896
rect 10428 18856 10692 18884
rect 10428 18828 10456 18856
rect 10686 18844 10692 18856
rect 10744 18844 10750 18896
rect 10962 18844 10968 18896
rect 11020 18884 11026 18896
rect 12084 18884 12112 18924
rect 12250 18912 12256 18964
rect 12308 18952 12314 18964
rect 15286 18952 15292 18964
rect 12308 18924 15292 18952
rect 12308 18912 12314 18924
rect 15286 18912 15292 18924
rect 15344 18912 15350 18964
rect 16853 18955 16911 18961
rect 16853 18921 16865 18955
rect 16899 18921 16911 18955
rect 16853 18915 16911 18921
rect 15304 18884 15332 18912
rect 11020 18856 12020 18884
rect 12084 18856 14688 18884
rect 15304 18856 16528 18884
rect 11020 18844 11026 18856
rect 8754 18816 8760 18828
rect 7944 18788 8760 18816
rect 7837 18779 7895 18785
rect 7374 18748 7380 18760
rect 6012 18720 6224 18748
rect 6472 18720 7380 18748
rect 5905 18711 5963 18717
rect 3145 18683 3203 18689
rect 3145 18649 3157 18683
rect 3191 18680 3203 18683
rect 3234 18680 3240 18692
rect 3191 18652 3240 18680
rect 3191 18649 3203 18652
rect 3145 18643 3203 18649
rect 3234 18640 3240 18652
rect 3292 18640 3298 18692
rect 4433 18683 4491 18689
rect 4433 18649 4445 18683
rect 4479 18680 4491 18683
rect 4890 18680 4896 18692
rect 4479 18652 4896 18680
rect 4479 18649 4491 18652
rect 4433 18643 4491 18649
rect 4890 18640 4896 18652
rect 4948 18640 4954 18692
rect 6196 18680 6224 18720
rect 7374 18708 7380 18720
rect 7432 18708 7438 18760
rect 6822 18680 6828 18692
rect 6196 18652 6828 18680
rect 6822 18640 6828 18652
rect 6880 18640 6886 18692
rect 6914 18640 6920 18692
rect 6972 18680 6978 18692
rect 7101 18683 7159 18689
rect 7101 18680 7113 18683
rect 6972 18652 7113 18680
rect 6972 18640 6978 18652
rect 7101 18649 7113 18652
rect 7147 18649 7159 18683
rect 7484 18680 7512 18779
rect 7558 18708 7564 18760
rect 7616 18748 7622 18760
rect 7852 18748 7880 18779
rect 8754 18776 8760 18788
rect 8812 18816 8818 18828
rect 8849 18819 8907 18825
rect 8849 18816 8861 18819
rect 8812 18788 8861 18816
rect 8812 18776 8818 18788
rect 8849 18785 8861 18788
rect 8895 18785 8907 18819
rect 8849 18779 8907 18785
rect 9582 18776 9588 18828
rect 9640 18776 9646 18828
rect 10410 18776 10416 18828
rect 10468 18776 10474 18828
rect 10594 18776 10600 18828
rect 10652 18776 10658 18828
rect 11054 18776 11060 18828
rect 11112 18816 11118 18828
rect 11992 18825 12020 18856
rect 11425 18819 11483 18825
rect 11425 18816 11437 18819
rect 11112 18788 11437 18816
rect 11112 18776 11118 18788
rect 11425 18785 11437 18788
rect 11471 18785 11483 18819
rect 11425 18779 11483 18785
rect 11977 18819 12035 18825
rect 11977 18785 11989 18819
rect 12023 18785 12035 18819
rect 11977 18779 12035 18785
rect 12158 18776 12164 18828
rect 12216 18776 12222 18828
rect 12710 18776 12716 18828
rect 12768 18776 12774 18828
rect 12986 18776 12992 18828
rect 13044 18776 13050 18828
rect 13143 18819 13201 18825
rect 13143 18785 13155 18819
rect 13189 18816 13201 18819
rect 13354 18816 13360 18828
rect 13189 18788 13360 18816
rect 13189 18785 13201 18788
rect 13143 18779 13201 18785
rect 13354 18776 13360 18788
rect 13412 18776 13418 18828
rect 14660 18825 14688 18856
rect 14645 18819 14703 18825
rect 14645 18785 14657 18819
rect 14691 18816 14703 18819
rect 15746 18816 15752 18828
rect 14691 18788 15752 18816
rect 14691 18785 14703 18788
rect 14645 18779 14703 18785
rect 15746 18776 15752 18788
rect 15804 18776 15810 18828
rect 16500 18825 16528 18856
rect 16485 18819 16543 18825
rect 16485 18785 16497 18819
rect 16531 18785 16543 18819
rect 16868 18816 16896 18915
rect 17310 18912 17316 18964
rect 17368 18952 17374 18964
rect 17681 18955 17739 18961
rect 17681 18952 17693 18955
rect 17368 18924 17693 18952
rect 17368 18912 17374 18924
rect 17681 18921 17693 18924
rect 17727 18952 17739 18955
rect 17954 18952 17960 18964
rect 17727 18924 17960 18952
rect 17727 18921 17739 18924
rect 17681 18915 17739 18921
rect 17954 18912 17960 18924
rect 18012 18912 18018 18964
rect 18414 18912 18420 18964
rect 18472 18912 18478 18964
rect 20346 18912 20352 18964
rect 20404 18952 20410 18964
rect 20625 18955 20683 18961
rect 20625 18952 20637 18955
rect 20404 18924 20637 18952
rect 20404 18912 20410 18924
rect 20625 18921 20637 18924
rect 20671 18952 20683 18955
rect 21450 18952 21456 18964
rect 20671 18924 21456 18952
rect 20671 18921 20683 18924
rect 20625 18915 20683 18921
rect 21450 18912 21456 18924
rect 21508 18912 21514 18964
rect 17770 18844 17776 18896
rect 17828 18884 17834 18896
rect 17865 18887 17923 18893
rect 17865 18884 17877 18887
rect 17828 18856 17877 18884
rect 17828 18844 17834 18856
rect 17865 18853 17877 18856
rect 17911 18853 17923 18887
rect 17865 18847 17923 18853
rect 19144 18887 19202 18893
rect 19144 18853 19156 18887
rect 19190 18884 19202 18887
rect 19242 18884 19248 18896
rect 19190 18856 19248 18884
rect 19190 18853 19202 18856
rect 19144 18847 19202 18853
rect 19242 18844 19248 18856
rect 19300 18844 19306 18896
rect 21634 18844 21640 18896
rect 21692 18884 21698 18896
rect 22382 18887 22440 18893
rect 22382 18884 22394 18887
rect 21692 18856 22394 18884
rect 21692 18844 21698 18856
rect 22382 18853 22394 18856
rect 22428 18853 22440 18887
rect 22382 18847 22440 18853
rect 17218 18816 17224 18828
rect 16868 18788 17224 18816
rect 16485 18779 16543 18785
rect 8478 18748 8484 18760
rect 7616 18720 7880 18748
rect 8036 18720 8484 18748
rect 7616 18708 7622 18720
rect 8036 18680 8064 18720
rect 8478 18708 8484 18720
rect 8536 18708 8542 18760
rect 11238 18708 11244 18760
rect 11296 18708 11302 18760
rect 11609 18751 11667 18757
rect 11609 18717 11621 18751
rect 11655 18748 11667 18751
rect 12437 18751 12495 18757
rect 12437 18748 12449 18751
rect 11655 18720 12449 18748
rect 11655 18717 11667 18720
rect 11609 18711 11667 18717
rect 12437 18717 12449 18720
rect 12483 18748 12495 18751
rect 12526 18748 12532 18760
rect 12483 18720 12532 18748
rect 12483 18717 12495 18720
rect 12437 18711 12495 18717
rect 12526 18708 12532 18720
rect 12584 18748 12590 18760
rect 13262 18748 13268 18760
rect 12584 18720 13268 18748
rect 12584 18708 12590 18720
rect 13262 18708 13268 18720
rect 13320 18708 13326 18760
rect 14550 18708 14556 18760
rect 14608 18708 14614 18760
rect 16390 18708 16396 18760
rect 16448 18708 16454 18760
rect 16500 18748 16528 18779
rect 17218 18776 17224 18788
rect 17276 18776 17282 18828
rect 17402 18776 17408 18828
rect 17460 18776 17466 18828
rect 17586 18776 17592 18828
rect 17644 18776 17650 18828
rect 18046 18776 18052 18828
rect 18104 18776 18110 18828
rect 18233 18819 18291 18825
rect 18233 18785 18245 18819
rect 18279 18816 18291 18819
rect 18325 18819 18383 18825
rect 18325 18816 18337 18819
rect 18279 18788 18337 18816
rect 18279 18785 18291 18788
rect 18233 18779 18291 18785
rect 18325 18785 18337 18788
rect 18371 18785 18383 18819
rect 18509 18819 18567 18825
rect 18509 18816 18521 18819
rect 18325 18779 18383 18785
rect 18432 18788 18521 18816
rect 17126 18748 17132 18760
rect 16500 18720 17132 18748
rect 17126 18708 17132 18720
rect 17184 18708 17190 18760
rect 18248 18748 18276 18779
rect 17880 18720 18276 18748
rect 9490 18680 9496 18692
rect 7484 18652 8064 18680
rect 8128 18652 9496 18680
rect 7101 18643 7159 18649
rect 3510 18572 3516 18624
rect 3568 18612 3574 18624
rect 3605 18615 3663 18621
rect 3605 18612 3617 18615
rect 3568 18584 3617 18612
rect 3568 18572 3574 18584
rect 3605 18581 3617 18584
rect 3651 18581 3663 18615
rect 3605 18575 3663 18581
rect 3973 18615 4031 18621
rect 3973 18581 3985 18615
rect 4019 18612 4031 18615
rect 4062 18612 4068 18624
rect 4019 18584 4068 18612
rect 4019 18581 4031 18584
rect 3973 18575 4031 18581
rect 4062 18572 4068 18584
rect 4120 18572 4126 18624
rect 7009 18615 7067 18621
rect 7009 18581 7021 18615
rect 7055 18612 7067 18615
rect 8128 18612 8156 18652
rect 9490 18640 9496 18652
rect 9548 18640 9554 18692
rect 13357 18683 13415 18689
rect 13357 18649 13369 18683
rect 13403 18680 13415 18683
rect 13906 18680 13912 18692
rect 13403 18652 13912 18680
rect 13403 18649 13415 18652
rect 13357 18643 13415 18649
rect 13906 18640 13912 18652
rect 13964 18640 13970 18692
rect 17880 18689 17908 18720
rect 17865 18683 17923 18689
rect 17865 18649 17877 18683
rect 17911 18649 17923 18683
rect 18432 18680 18460 18788
rect 18509 18785 18521 18788
rect 18555 18785 18567 18819
rect 18509 18779 18567 18785
rect 19610 18776 19616 18828
rect 19668 18816 19674 18828
rect 20809 18819 20867 18825
rect 20809 18816 20821 18819
rect 19668 18788 20821 18816
rect 19668 18776 19674 18788
rect 20809 18785 20821 18788
rect 20855 18785 20867 18819
rect 20809 18779 20867 18785
rect 20993 18819 21051 18825
rect 20993 18785 21005 18819
rect 21039 18816 21051 18819
rect 21266 18816 21272 18828
rect 21039 18788 21272 18816
rect 21039 18785 21051 18788
rect 20993 18779 21051 18785
rect 21266 18776 21272 18788
rect 21324 18776 21330 18828
rect 22925 18819 22983 18825
rect 22925 18816 22937 18819
rect 22664 18788 22937 18816
rect 22664 18760 22692 18788
rect 22925 18785 22937 18788
rect 22971 18785 22983 18819
rect 22925 18779 22983 18785
rect 18874 18708 18880 18760
rect 18932 18708 18938 18760
rect 20898 18708 20904 18760
rect 20956 18748 20962 18760
rect 21085 18751 21143 18757
rect 21085 18748 21097 18751
rect 20956 18720 21097 18748
rect 20956 18708 20962 18720
rect 21085 18717 21097 18720
rect 21131 18717 21143 18751
rect 21085 18711 21143 18717
rect 22646 18708 22652 18760
rect 22704 18708 22710 18760
rect 17865 18643 17923 18649
rect 18156 18652 18460 18680
rect 7055 18584 8156 18612
rect 7055 18581 7067 18584
rect 7009 18575 7067 18581
rect 8202 18572 8208 18624
rect 8260 18572 8266 18624
rect 8294 18572 8300 18624
rect 8352 18572 8358 18624
rect 10042 18572 10048 18624
rect 10100 18612 10106 18624
rect 10413 18615 10471 18621
rect 10413 18612 10425 18615
rect 10100 18584 10425 18612
rect 10100 18572 10106 18584
rect 10413 18581 10425 18584
rect 10459 18581 10471 18615
rect 10413 18575 10471 18581
rect 12345 18615 12403 18621
rect 12345 18581 12357 18615
rect 12391 18612 12403 18615
rect 12529 18615 12587 18621
rect 12529 18612 12541 18615
rect 12391 18584 12541 18612
rect 12391 18581 12403 18584
rect 12345 18575 12403 18581
rect 12529 18581 12541 18584
rect 12575 18612 12587 18615
rect 12618 18612 12624 18624
rect 12575 18584 12624 18612
rect 12575 18581 12587 18584
rect 12529 18575 12587 18581
rect 12618 18572 12624 18584
rect 12676 18572 12682 18624
rect 12894 18572 12900 18624
rect 12952 18572 12958 18624
rect 15010 18572 15016 18624
rect 15068 18572 15074 18624
rect 17405 18615 17463 18621
rect 17405 18581 17417 18615
rect 17451 18612 17463 18615
rect 17770 18612 17776 18624
rect 17451 18584 17776 18612
rect 17451 18581 17463 18584
rect 17405 18575 17463 18581
rect 17770 18572 17776 18584
rect 17828 18612 17834 18624
rect 18156 18612 18184 18652
rect 17828 18584 18184 18612
rect 18233 18615 18291 18621
rect 17828 18572 17834 18584
rect 18233 18581 18245 18615
rect 18279 18612 18291 18615
rect 18414 18612 18420 18624
rect 18279 18584 18420 18612
rect 18279 18581 18291 18584
rect 18233 18575 18291 18581
rect 18414 18572 18420 18584
rect 18472 18572 18478 18624
rect 20070 18572 20076 18624
rect 20128 18612 20134 18624
rect 20257 18615 20315 18621
rect 20257 18612 20269 18615
rect 20128 18584 20269 18612
rect 20128 18572 20134 18584
rect 20257 18581 20269 18584
rect 20303 18581 20315 18615
rect 20257 18575 20315 18581
rect 21082 18572 21088 18624
rect 21140 18612 21146 18624
rect 21269 18615 21327 18621
rect 21269 18612 21281 18615
rect 21140 18584 21281 18612
rect 21140 18572 21146 18584
rect 21269 18581 21281 18584
rect 21315 18581 21327 18615
rect 21269 18575 21327 18581
rect 21634 18572 21640 18624
rect 21692 18612 21698 18624
rect 22278 18612 22284 18624
rect 21692 18584 22284 18612
rect 21692 18572 21698 18584
rect 22278 18572 22284 18584
rect 22336 18612 22342 18624
rect 22833 18615 22891 18621
rect 22833 18612 22845 18615
rect 22336 18584 22845 18612
rect 22336 18572 22342 18584
rect 22833 18581 22845 18584
rect 22879 18581 22891 18615
rect 22833 18575 22891 18581
rect 552 18522 23368 18544
rect 552 18470 3662 18522
rect 3714 18470 3726 18522
rect 3778 18470 3790 18522
rect 3842 18470 3854 18522
rect 3906 18470 3918 18522
rect 3970 18470 23368 18522
rect 552 18448 23368 18470
rect 5445 18411 5503 18417
rect 5445 18377 5457 18411
rect 5491 18408 5503 18411
rect 6270 18408 6276 18420
rect 5491 18380 6276 18408
rect 5491 18377 5503 18380
rect 5445 18371 5503 18377
rect 6270 18368 6276 18380
rect 6328 18368 6334 18420
rect 12618 18368 12624 18420
rect 12676 18408 12682 18420
rect 12676 18380 13032 18408
rect 12676 18368 12682 18380
rect 9582 18300 9588 18352
rect 9640 18300 9646 18352
rect 10042 18300 10048 18352
rect 10100 18340 10106 18352
rect 11885 18343 11943 18349
rect 10100 18312 11560 18340
rect 10100 18300 10106 18312
rect 3326 18232 3332 18284
rect 3384 18272 3390 18284
rect 3421 18275 3479 18281
rect 3421 18272 3433 18275
rect 3384 18244 3433 18272
rect 3384 18232 3390 18244
rect 3421 18241 3433 18244
rect 3467 18241 3479 18275
rect 3421 18235 3479 18241
rect 3881 18275 3939 18281
rect 3881 18241 3893 18275
rect 3927 18272 3939 18275
rect 4246 18272 4252 18284
rect 3927 18244 4252 18272
rect 3927 18241 3939 18244
rect 3881 18235 3939 18241
rect 4246 18232 4252 18244
rect 4304 18232 4310 18284
rect 7374 18232 7380 18284
rect 7432 18272 7438 18284
rect 9401 18275 9459 18281
rect 7432 18244 7604 18272
rect 7432 18232 7438 18244
rect 3513 18207 3571 18213
rect 3513 18173 3525 18207
rect 3559 18204 3571 18207
rect 4338 18204 4344 18216
rect 3559 18176 4344 18204
rect 3559 18173 3571 18176
rect 3513 18167 3571 18173
rect 4338 18164 4344 18176
rect 4396 18204 4402 18216
rect 4890 18204 4896 18216
rect 4396 18176 4896 18204
rect 4396 18164 4402 18176
rect 4890 18164 4896 18176
rect 4948 18164 4954 18216
rect 5258 18164 5264 18216
rect 5316 18164 5322 18216
rect 7282 18164 7288 18216
rect 7340 18164 7346 18216
rect 7466 18164 7472 18216
rect 7524 18164 7530 18216
rect 7576 18213 7604 18244
rect 9401 18241 9413 18275
rect 9447 18272 9459 18275
rect 9600 18272 9628 18300
rect 9447 18244 9628 18272
rect 9447 18241 9459 18244
rect 9401 18235 9459 18241
rect 9950 18232 9956 18284
rect 10008 18272 10014 18284
rect 10505 18275 10563 18281
rect 10505 18272 10517 18275
rect 10008 18244 10517 18272
rect 10008 18232 10014 18244
rect 10505 18241 10517 18244
rect 10551 18272 10563 18275
rect 11425 18275 11483 18281
rect 11425 18272 11437 18275
rect 10551 18244 11437 18272
rect 10551 18241 10563 18244
rect 10505 18235 10563 18241
rect 11425 18241 11437 18244
rect 11471 18241 11483 18275
rect 11425 18235 11483 18241
rect 7561 18207 7619 18213
rect 7561 18173 7573 18207
rect 7607 18173 7619 18207
rect 7561 18167 7619 18173
rect 7745 18207 7803 18213
rect 7745 18173 7757 18207
rect 7791 18204 7803 18207
rect 8386 18204 8392 18216
rect 7791 18176 8392 18204
rect 7791 18173 7803 18176
rect 7745 18167 7803 18173
rect 8386 18164 8392 18176
rect 8444 18164 8450 18216
rect 8754 18164 8760 18216
rect 8812 18164 8818 18216
rect 9585 18207 9643 18213
rect 9585 18173 9597 18207
rect 9631 18173 9643 18207
rect 9585 18167 9643 18173
rect 5074 18096 5080 18148
rect 5132 18096 5138 18148
rect 8665 18139 8723 18145
rect 8665 18105 8677 18139
rect 8711 18136 8723 18139
rect 9030 18136 9036 18148
rect 8711 18108 9036 18136
rect 8711 18105 8723 18108
rect 8665 18099 8723 18105
rect 9030 18096 9036 18108
rect 9088 18136 9094 18148
rect 9600 18136 9628 18167
rect 10042 18164 10048 18216
rect 10100 18164 10106 18216
rect 10410 18164 10416 18216
rect 10468 18204 10474 18216
rect 10597 18207 10655 18213
rect 10597 18204 10609 18207
rect 10468 18176 10609 18204
rect 10468 18164 10474 18176
rect 10597 18173 10609 18176
rect 10643 18173 10655 18207
rect 10597 18167 10655 18173
rect 10686 18164 10692 18216
rect 10744 18204 10750 18216
rect 10781 18207 10839 18213
rect 10781 18204 10793 18207
rect 10744 18176 10793 18204
rect 10744 18164 10750 18176
rect 10781 18173 10793 18176
rect 10827 18173 10839 18207
rect 10781 18167 10839 18173
rect 11146 18164 11152 18216
rect 11204 18164 11210 18216
rect 11532 18213 11560 18312
rect 11885 18309 11897 18343
rect 11931 18309 11943 18343
rect 11885 18303 11943 18309
rect 11900 18272 11928 18303
rect 12434 18300 12440 18352
rect 12492 18340 12498 18352
rect 13004 18349 13032 18380
rect 19702 18368 19708 18420
rect 19760 18368 19766 18420
rect 20990 18368 20996 18420
rect 21048 18368 21054 18420
rect 21174 18368 21180 18420
rect 21232 18408 21238 18420
rect 22278 18408 22284 18420
rect 21232 18380 22284 18408
rect 21232 18368 21238 18380
rect 22278 18368 22284 18380
rect 22336 18408 22342 18420
rect 23017 18411 23075 18417
rect 23017 18408 23029 18411
rect 22336 18380 23029 18408
rect 22336 18368 22342 18380
rect 23017 18377 23029 18380
rect 23063 18377 23075 18411
rect 23017 18371 23075 18377
rect 12897 18343 12955 18349
rect 12897 18340 12909 18343
rect 12492 18312 12909 18340
rect 12492 18300 12498 18312
rect 12897 18309 12909 18312
rect 12943 18309 12955 18343
rect 12897 18303 12955 18309
rect 12989 18343 13047 18349
rect 12989 18309 13001 18343
rect 13035 18309 13047 18343
rect 12989 18303 13047 18309
rect 13078 18300 13084 18352
rect 13136 18340 13142 18352
rect 13817 18343 13875 18349
rect 13136 18312 13768 18340
rect 13136 18300 13142 18312
rect 12710 18272 12716 18284
rect 11900 18244 12716 18272
rect 12710 18232 12716 18244
rect 12768 18272 12774 18284
rect 12805 18275 12863 18281
rect 12805 18272 12817 18275
rect 12768 18244 12817 18272
rect 12768 18232 12774 18244
rect 12805 18241 12817 18244
rect 12851 18272 12863 18275
rect 13173 18275 13231 18281
rect 12851 18244 13032 18272
rect 12851 18241 12863 18244
rect 12805 18235 12863 18241
rect 11517 18207 11575 18213
rect 11517 18173 11529 18207
rect 11563 18173 11575 18207
rect 11517 18167 11575 18173
rect 12526 18164 12532 18216
rect 12584 18164 12590 18216
rect 12897 18207 12955 18213
rect 12897 18173 12909 18207
rect 12943 18206 12955 18207
rect 13004 18206 13032 18244
rect 13173 18241 13185 18275
rect 13219 18272 13231 18275
rect 13262 18272 13268 18284
rect 13219 18244 13268 18272
rect 13219 18241 13231 18244
rect 13173 18235 13231 18241
rect 13262 18232 13268 18244
rect 13320 18232 13326 18284
rect 13740 18272 13768 18312
rect 13817 18309 13829 18343
rect 13863 18340 13875 18343
rect 14918 18340 14924 18352
rect 13863 18312 14924 18340
rect 13863 18309 13875 18312
rect 13817 18303 13875 18309
rect 14918 18300 14924 18312
rect 14976 18300 14982 18352
rect 15286 18300 15292 18352
rect 15344 18340 15350 18352
rect 16485 18343 16543 18349
rect 15344 18312 16344 18340
rect 15344 18300 15350 18312
rect 13740 18244 14136 18272
rect 14108 18213 14136 18244
rect 15010 18232 15016 18284
rect 15068 18272 15074 18284
rect 15381 18275 15439 18281
rect 15381 18272 15393 18275
rect 15068 18244 15393 18272
rect 15068 18232 15074 18244
rect 15381 18241 15393 18244
rect 15427 18272 15439 18275
rect 15427 18244 16252 18272
rect 15427 18241 15439 18244
rect 15381 18235 15439 18241
rect 12943 18178 13032 18206
rect 13541 18207 13599 18213
rect 13541 18204 13553 18207
rect 12943 18173 12955 18178
rect 12897 18167 12955 18173
rect 13188 18176 13553 18204
rect 9088 18108 9628 18136
rect 10321 18139 10379 18145
rect 9088 18096 9094 18108
rect 10321 18105 10333 18139
rect 10367 18136 10379 18139
rect 11054 18136 11060 18148
rect 10367 18108 11060 18136
rect 10367 18105 10379 18108
rect 10321 18099 10379 18105
rect 11054 18096 11060 18108
rect 11112 18136 11118 18148
rect 12250 18136 12256 18148
rect 11112 18108 12256 18136
rect 11112 18096 11118 18108
rect 12250 18096 12256 18108
rect 12308 18096 12314 18148
rect 12805 18139 12863 18145
rect 12805 18105 12817 18139
rect 12851 18105 12863 18139
rect 13188 18136 13216 18176
rect 13541 18173 13553 18176
rect 13587 18173 13599 18207
rect 13541 18167 13599 18173
rect 13909 18207 13967 18213
rect 13909 18173 13921 18207
rect 13955 18173 13967 18207
rect 13909 18167 13967 18173
rect 14093 18207 14151 18213
rect 14093 18173 14105 18207
rect 14139 18173 14151 18207
rect 14093 18167 14151 18173
rect 12805 18099 12863 18105
rect 13004 18108 13216 18136
rect 7374 18028 7380 18080
rect 7432 18028 7438 18080
rect 7742 18028 7748 18080
rect 7800 18028 7806 18080
rect 11241 18071 11299 18077
rect 11241 18037 11253 18071
rect 11287 18068 11299 18071
rect 12158 18068 12164 18080
rect 11287 18040 12164 18068
rect 11287 18037 11299 18040
rect 11241 18031 11299 18037
rect 12158 18028 12164 18040
rect 12216 18028 12222 18080
rect 12820 18068 12848 18099
rect 13004 18068 13032 18108
rect 13446 18096 13452 18148
rect 13504 18136 13510 18148
rect 13817 18139 13875 18145
rect 13817 18136 13829 18139
rect 13504 18108 13829 18136
rect 13504 18096 13510 18108
rect 13817 18105 13829 18108
rect 13863 18136 13875 18139
rect 13924 18136 13952 18167
rect 15286 18164 15292 18216
rect 15344 18164 15350 18216
rect 15746 18164 15752 18216
rect 15804 18164 15810 18216
rect 16224 18213 16252 18244
rect 16316 18213 16344 18312
rect 16485 18309 16497 18343
rect 16531 18309 16543 18343
rect 16485 18303 16543 18309
rect 15933 18207 15991 18213
rect 15933 18173 15945 18207
rect 15979 18173 15991 18207
rect 15933 18167 15991 18173
rect 16209 18207 16267 18213
rect 16209 18173 16221 18207
rect 16255 18173 16267 18207
rect 16209 18167 16267 18173
rect 16301 18207 16359 18213
rect 16301 18173 16313 18207
rect 16347 18173 16359 18207
rect 16500 18204 16528 18303
rect 17218 18232 17224 18284
rect 17276 18232 17282 18284
rect 20806 18272 20812 18284
rect 19904 18244 20812 18272
rect 19904 18216 19932 18244
rect 20806 18232 20812 18244
rect 20864 18272 20870 18284
rect 20864 18244 20944 18272
rect 20864 18232 20870 18244
rect 17402 18204 17408 18216
rect 16500 18176 17408 18204
rect 16301 18167 16359 18173
rect 13863 18108 13952 18136
rect 13863 18105 13875 18108
rect 13817 18099 13875 18105
rect 14550 18096 14556 18148
rect 14608 18136 14614 18148
rect 15948 18136 15976 18167
rect 17402 18164 17408 18176
rect 17460 18164 17466 18216
rect 19886 18164 19892 18216
rect 19944 18164 19950 18216
rect 20070 18164 20076 18216
rect 20128 18164 20134 18216
rect 20916 18213 20944 18244
rect 21358 18232 21364 18284
rect 21416 18272 21422 18284
rect 21416 18244 21772 18272
rect 21416 18232 21422 18244
rect 20901 18207 20959 18213
rect 20901 18173 20913 18207
rect 20947 18173 20959 18207
rect 20901 18167 20959 18173
rect 21634 18164 21640 18216
rect 21692 18164 21698 18216
rect 21744 18204 21772 18244
rect 21893 18207 21951 18213
rect 21893 18204 21905 18207
rect 21744 18176 21905 18204
rect 21893 18173 21905 18176
rect 21939 18173 21951 18207
rect 21893 18167 21951 18173
rect 14608 18108 15976 18136
rect 16117 18139 16175 18145
rect 14608 18096 14614 18108
rect 16117 18105 16129 18139
rect 16163 18136 16175 18139
rect 16485 18139 16543 18145
rect 16485 18136 16497 18139
rect 16163 18108 16497 18136
rect 16163 18105 16175 18108
rect 16117 18099 16175 18105
rect 16485 18105 16497 18108
rect 16531 18105 16543 18139
rect 16485 18099 16543 18105
rect 18874 18096 18880 18148
rect 18932 18136 18938 18148
rect 21652 18136 21680 18164
rect 18932 18108 21680 18136
rect 18932 18096 18938 18108
rect 12820 18040 13032 18068
rect 13633 18071 13691 18077
rect 13633 18037 13645 18071
rect 13679 18068 13691 18071
rect 13906 18068 13912 18080
rect 13679 18040 13912 18068
rect 13679 18037 13691 18040
rect 13633 18031 13691 18037
rect 13906 18028 13912 18040
rect 13964 18028 13970 18080
rect 13998 18028 14004 18080
rect 14056 18028 14062 18080
rect 15654 18028 15660 18080
rect 15712 18028 15718 18080
rect 17589 18071 17647 18077
rect 17589 18037 17601 18071
rect 17635 18068 17647 18071
rect 17678 18068 17684 18080
rect 17635 18040 17684 18068
rect 17635 18037 17647 18040
rect 17589 18031 17647 18037
rect 17678 18028 17684 18040
rect 17736 18028 17742 18080
rect 552 17978 23368 18000
rect 552 17926 4322 17978
rect 4374 17926 4386 17978
rect 4438 17926 4450 17978
rect 4502 17926 4514 17978
rect 4566 17926 4578 17978
rect 4630 17926 23368 17978
rect 552 17904 23368 17926
rect 4249 17867 4307 17873
rect 4249 17833 4261 17867
rect 4295 17864 4307 17867
rect 5074 17864 5080 17876
rect 4295 17836 5080 17864
rect 4295 17833 4307 17836
rect 4249 17827 4307 17833
rect 5074 17824 5080 17836
rect 5132 17824 5138 17876
rect 10413 17867 10471 17873
rect 10413 17833 10425 17867
rect 10459 17864 10471 17867
rect 11146 17864 11152 17876
rect 10459 17836 11152 17864
rect 10459 17833 10471 17836
rect 10413 17827 10471 17833
rect 11146 17824 11152 17836
rect 11204 17824 11210 17876
rect 14093 17867 14151 17873
rect 14093 17833 14105 17867
rect 14139 17864 14151 17867
rect 15286 17864 15292 17876
rect 14139 17836 15292 17864
rect 14139 17833 14151 17836
rect 14093 17827 14151 17833
rect 15286 17824 15292 17836
rect 15344 17824 15350 17876
rect 2774 17756 2780 17808
rect 2832 17796 2838 17808
rect 3418 17796 3424 17808
rect 2832 17768 3424 17796
rect 2832 17756 2838 17768
rect 3418 17756 3424 17768
rect 3476 17796 3482 17808
rect 3476 17768 3832 17796
rect 3476 17756 3482 17768
rect 3326 17688 3332 17740
rect 3384 17728 3390 17740
rect 3804 17737 3832 17768
rect 9490 17756 9496 17808
rect 9548 17796 9554 17808
rect 13446 17796 13452 17808
rect 9548 17768 10272 17796
rect 9548 17756 9554 17768
rect 3605 17731 3663 17737
rect 3605 17728 3617 17731
rect 3384 17700 3617 17728
rect 3384 17688 3390 17700
rect 3605 17697 3617 17700
rect 3651 17697 3663 17731
rect 3605 17691 3663 17697
rect 3789 17731 3847 17737
rect 3789 17697 3801 17731
rect 3835 17697 3847 17731
rect 3789 17691 3847 17697
rect 4065 17731 4123 17737
rect 4065 17697 4077 17731
rect 4111 17697 4123 17731
rect 4065 17691 4123 17697
rect 3142 17620 3148 17672
rect 3200 17660 3206 17672
rect 4080 17660 4108 17691
rect 9582 17688 9588 17740
rect 9640 17728 9646 17740
rect 10244 17737 10272 17768
rect 13096 17768 13452 17796
rect 10045 17731 10103 17737
rect 10045 17728 10057 17731
rect 9640 17700 10057 17728
rect 9640 17688 9646 17700
rect 10045 17697 10057 17700
rect 10091 17697 10103 17731
rect 10045 17691 10103 17697
rect 10229 17731 10287 17737
rect 10229 17697 10241 17731
rect 10275 17697 10287 17731
rect 10229 17691 10287 17697
rect 12434 17688 12440 17740
rect 12492 17728 12498 17740
rect 13096 17737 13124 17768
rect 13446 17756 13452 17768
rect 13504 17756 13510 17808
rect 13906 17756 13912 17808
rect 13964 17796 13970 17808
rect 21821 17799 21879 17805
rect 13964 17768 14504 17796
rect 13964 17756 13970 17768
rect 13081 17731 13139 17737
rect 13081 17728 13093 17731
rect 12492 17700 13093 17728
rect 12492 17688 12498 17700
rect 13081 17697 13093 17700
rect 13127 17697 13139 17731
rect 13081 17691 13139 17697
rect 13170 17688 13176 17740
rect 13228 17688 13234 17740
rect 13725 17731 13783 17737
rect 13725 17697 13737 17731
rect 13771 17728 13783 17731
rect 13998 17728 14004 17740
rect 13771 17700 14004 17728
rect 13771 17697 13783 17700
rect 13725 17691 13783 17697
rect 13998 17688 14004 17700
rect 14056 17688 14062 17740
rect 14476 17737 14504 17768
rect 21821 17765 21833 17799
rect 21867 17796 21879 17799
rect 22094 17796 22100 17808
rect 21867 17768 22100 17796
rect 21867 17765 21879 17768
rect 21821 17759 21879 17765
rect 22094 17756 22100 17768
rect 22152 17796 22158 17808
rect 22830 17796 22836 17808
rect 22152 17768 22836 17796
rect 22152 17756 22158 17768
rect 22830 17756 22836 17768
rect 22888 17756 22894 17808
rect 14461 17731 14519 17737
rect 14461 17697 14473 17731
rect 14507 17697 14519 17731
rect 14461 17691 14519 17697
rect 17678 17688 17684 17740
rect 17736 17688 17742 17740
rect 17770 17688 17776 17740
rect 17828 17728 17834 17740
rect 17865 17731 17923 17737
rect 17865 17728 17877 17731
rect 17828 17700 17877 17728
rect 17828 17688 17834 17700
rect 17865 17697 17877 17700
rect 17911 17697 17923 17731
rect 17865 17691 17923 17697
rect 21634 17688 21640 17740
rect 21692 17688 21698 17740
rect 21913 17731 21971 17737
rect 21913 17697 21925 17731
rect 21959 17728 21971 17731
rect 22002 17728 22008 17740
rect 21959 17700 22008 17728
rect 21959 17697 21971 17700
rect 21913 17691 21971 17697
rect 22002 17688 22008 17700
rect 22060 17688 22066 17740
rect 3200 17632 4108 17660
rect 3200 17620 3206 17632
rect 9490 17620 9496 17672
rect 9548 17620 9554 17672
rect 9950 17620 9956 17672
rect 10008 17620 10014 17672
rect 13633 17663 13691 17669
rect 13633 17629 13645 17663
rect 13679 17629 13691 17663
rect 13633 17623 13691 17629
rect 13648 17592 13676 17623
rect 13906 17620 13912 17672
rect 13964 17660 13970 17672
rect 14185 17663 14243 17669
rect 14185 17660 14197 17663
rect 13964 17632 14197 17660
rect 13964 17620 13970 17632
rect 14185 17629 14197 17632
rect 14231 17629 14243 17663
rect 14185 17623 14243 17629
rect 14645 17595 14703 17601
rect 14645 17592 14657 17595
rect 13648 17564 14657 17592
rect 14645 17561 14657 17564
rect 14691 17561 14703 17595
rect 14645 17555 14703 17561
rect 12894 17484 12900 17536
rect 12952 17524 12958 17536
rect 13081 17527 13139 17533
rect 13081 17524 13093 17527
rect 12952 17496 13093 17524
rect 12952 17484 12958 17496
rect 13081 17493 13093 17496
rect 13127 17493 13139 17527
rect 13081 17487 13139 17493
rect 13449 17527 13507 17533
rect 13449 17493 13461 17527
rect 13495 17524 13507 17527
rect 13998 17524 14004 17536
rect 13495 17496 14004 17524
rect 13495 17493 13507 17496
rect 13449 17487 13507 17493
rect 13998 17484 14004 17496
rect 14056 17484 14062 17536
rect 14274 17484 14280 17536
rect 14332 17484 14338 17536
rect 17681 17527 17739 17533
rect 17681 17493 17693 17527
rect 17727 17524 17739 17527
rect 17862 17524 17868 17536
rect 17727 17496 17868 17524
rect 17727 17493 17739 17496
rect 17681 17487 17739 17493
rect 17862 17484 17868 17496
rect 17920 17484 17926 17536
rect 21637 17527 21695 17533
rect 21637 17493 21649 17527
rect 21683 17524 21695 17527
rect 21726 17524 21732 17536
rect 21683 17496 21732 17524
rect 21683 17493 21695 17496
rect 21637 17487 21695 17493
rect 21726 17484 21732 17496
rect 21784 17484 21790 17536
rect 552 17434 23368 17456
rect 552 17382 3662 17434
rect 3714 17382 3726 17434
rect 3778 17382 3790 17434
rect 3842 17382 3854 17434
rect 3906 17382 3918 17434
rect 3970 17382 23368 17434
rect 552 17360 23368 17382
rect 3510 17280 3516 17332
rect 3568 17320 3574 17332
rect 3881 17323 3939 17329
rect 3881 17320 3893 17323
rect 3568 17292 3893 17320
rect 3568 17280 3574 17292
rect 3881 17289 3893 17292
rect 3927 17289 3939 17323
rect 3881 17283 3939 17289
rect 8849 17323 8907 17329
rect 8849 17289 8861 17323
rect 8895 17320 8907 17323
rect 9582 17320 9588 17332
rect 8895 17292 9588 17320
rect 8895 17289 8907 17292
rect 8849 17283 8907 17289
rect 9582 17280 9588 17292
rect 9640 17280 9646 17332
rect 9674 17280 9680 17332
rect 9732 17320 9738 17332
rect 14550 17320 14556 17332
rect 9732 17292 14556 17320
rect 9732 17280 9738 17292
rect 14550 17280 14556 17292
rect 14608 17280 14614 17332
rect 18414 17280 18420 17332
rect 18472 17320 18478 17332
rect 20714 17320 20720 17332
rect 18472 17292 19104 17320
rect 18472 17280 18478 17292
rect 14274 17252 14280 17264
rect 13648 17224 14280 17252
rect 7006 17144 7012 17196
rect 7064 17184 7070 17196
rect 8110 17184 8116 17196
rect 7064 17156 8116 17184
rect 7064 17144 7070 17156
rect 8110 17144 8116 17156
rect 8168 17184 8174 17196
rect 8481 17187 8539 17193
rect 8481 17184 8493 17187
rect 8168 17156 8493 17184
rect 8168 17144 8174 17156
rect 8481 17153 8493 17156
rect 8527 17153 8539 17187
rect 8481 17147 8539 17153
rect 13538 17144 13544 17196
rect 13596 17184 13602 17196
rect 13648 17193 13676 17224
rect 14274 17212 14280 17224
rect 14332 17212 14338 17264
rect 16758 17252 16764 17264
rect 15028 17224 16764 17252
rect 13633 17187 13691 17193
rect 13633 17184 13645 17187
rect 13596 17156 13645 17184
rect 13596 17144 13602 17156
rect 13633 17153 13645 17156
rect 13679 17153 13691 17187
rect 13633 17147 13691 17153
rect 14090 17144 14096 17196
rect 14148 17144 14154 17196
rect 5442 17076 5448 17128
rect 5500 17116 5506 17128
rect 5905 17119 5963 17125
rect 5905 17116 5917 17119
rect 5500 17088 5917 17116
rect 5500 17076 5506 17088
rect 5905 17085 5917 17088
rect 5951 17085 5963 17119
rect 5905 17079 5963 17085
rect 6086 17076 6092 17128
rect 6144 17076 6150 17128
rect 8573 17119 8631 17125
rect 8573 17085 8585 17119
rect 8619 17116 8631 17119
rect 8846 17116 8852 17128
rect 8619 17088 8852 17116
rect 8619 17085 8631 17088
rect 8573 17079 8631 17085
rect 8846 17076 8852 17088
rect 8904 17076 8910 17128
rect 13170 17076 13176 17128
rect 13228 17116 13234 17128
rect 13722 17116 13728 17128
rect 13228 17088 13728 17116
rect 13228 17076 13234 17088
rect 13722 17076 13728 17088
rect 13780 17076 13786 17128
rect 3326 17008 3332 17060
rect 3384 17048 3390 17060
rect 3602 17048 3608 17060
rect 3384 17020 3608 17048
rect 3384 17008 3390 17020
rect 3602 17008 3608 17020
rect 3660 17048 3666 17060
rect 3697 17051 3755 17057
rect 3697 17048 3709 17051
rect 3660 17020 3709 17048
rect 3660 17008 3666 17020
rect 3697 17017 3709 17020
rect 3743 17017 3755 17051
rect 3697 17011 3755 17017
rect 13630 17008 13636 17060
rect 13688 17048 13694 17060
rect 15028 17048 15056 17224
rect 16758 17212 16764 17224
rect 16816 17212 16822 17264
rect 19076 17261 19104 17292
rect 20364 17292 20720 17320
rect 18233 17255 18291 17261
rect 18233 17221 18245 17255
rect 18279 17252 18291 17255
rect 19061 17255 19119 17261
rect 18279 17224 19012 17252
rect 18279 17221 18291 17224
rect 18233 17215 18291 17221
rect 15654 17144 15660 17196
rect 15712 17144 15718 17196
rect 17770 17144 17776 17196
rect 17828 17184 17834 17196
rect 17828 17156 18184 17184
rect 17828 17144 17834 17156
rect 15841 17119 15899 17125
rect 15841 17116 15853 17119
rect 13688 17020 15056 17048
rect 15120 17088 15853 17116
rect 13688 17008 13694 17020
rect 15120 16992 15148 17088
rect 15841 17085 15853 17088
rect 15887 17085 15899 17119
rect 15841 17079 15899 17085
rect 17862 17076 17868 17128
rect 17920 17076 17926 17128
rect 18156 17125 18184 17156
rect 18414 17144 18420 17196
rect 18472 17144 18478 17196
rect 18984 17128 19012 17224
rect 19061 17221 19073 17255
rect 19107 17221 19119 17255
rect 19061 17215 19119 17221
rect 19610 17184 19616 17196
rect 19168 17156 19616 17184
rect 18049 17119 18107 17125
rect 18049 17085 18061 17119
rect 18095 17085 18107 17119
rect 18049 17079 18107 17085
rect 18141 17119 18199 17125
rect 18141 17085 18153 17119
rect 18187 17116 18199 17119
rect 18877 17119 18935 17125
rect 18877 17116 18889 17119
rect 18187 17088 18889 17116
rect 18187 17085 18199 17088
rect 18141 17079 18199 17085
rect 18877 17085 18889 17088
rect 18923 17085 18935 17119
rect 18877 17079 18935 17085
rect 18064 17048 18092 17079
rect 18966 17076 18972 17128
rect 19024 17076 19030 17128
rect 19058 17076 19064 17128
rect 19116 17116 19122 17128
rect 19168 17125 19196 17156
rect 19610 17144 19616 17156
rect 19668 17184 19674 17196
rect 19981 17187 20039 17193
rect 19981 17184 19993 17187
rect 19668 17156 19993 17184
rect 19668 17144 19674 17156
rect 19981 17153 19993 17156
rect 20027 17153 20039 17187
rect 19981 17147 20039 17153
rect 19153 17119 19211 17125
rect 19153 17116 19165 17119
rect 19116 17088 19165 17116
rect 19116 17076 19122 17088
rect 19153 17085 19165 17088
rect 19199 17085 19211 17119
rect 19153 17079 19211 17085
rect 19889 17119 19947 17125
rect 19889 17085 19901 17119
rect 19935 17085 19947 17119
rect 19889 17079 19947 17085
rect 20165 17119 20223 17125
rect 20165 17085 20177 17119
rect 20211 17116 20223 17119
rect 20364 17116 20392 17292
rect 20714 17280 20720 17292
rect 20772 17280 20778 17332
rect 22830 17280 22836 17332
rect 22888 17280 22894 17332
rect 20211 17088 20392 17116
rect 20211 17085 20223 17088
rect 20165 17079 20223 17085
rect 18322 17048 18328 17060
rect 18064 17020 18328 17048
rect 18322 17008 18328 17020
rect 18380 17008 18386 17060
rect 18417 17051 18475 17057
rect 18417 17017 18429 17051
rect 18463 17048 18475 17051
rect 18782 17048 18788 17060
rect 18463 17020 18788 17048
rect 18463 17017 18475 17020
rect 18417 17011 18475 17017
rect 18782 17008 18788 17020
rect 18840 17008 18846 17060
rect 3418 16940 3424 16992
rect 3476 16980 3482 16992
rect 3897 16983 3955 16989
rect 3897 16980 3909 16983
rect 3476 16952 3909 16980
rect 3476 16940 3482 16952
rect 3897 16949 3909 16952
rect 3943 16949 3955 16983
rect 3897 16943 3955 16949
rect 4062 16940 4068 16992
rect 4120 16940 4126 16992
rect 5997 16983 6055 16989
rect 5997 16949 6009 16983
rect 6043 16980 6055 16983
rect 7466 16980 7472 16992
rect 6043 16952 7472 16980
rect 6043 16949 6055 16952
rect 5997 16943 6055 16949
rect 7466 16940 7472 16952
rect 7524 16940 7530 16992
rect 11514 16940 11520 16992
rect 11572 16980 11578 16992
rect 15102 16980 15108 16992
rect 11572 16952 15108 16980
rect 11572 16940 11578 16952
rect 15102 16940 15108 16952
rect 15160 16940 15166 16992
rect 16022 16940 16028 16992
rect 16080 16940 16086 16992
rect 17954 16940 17960 16992
rect 18012 16940 18018 16992
rect 18690 16940 18696 16992
rect 18748 16940 18754 16992
rect 19904 16980 19932 17079
rect 20438 17076 20444 17128
rect 20496 17076 20502 17128
rect 22370 17076 22376 17128
rect 22428 17116 22434 17128
rect 22741 17119 22799 17125
rect 22741 17116 22753 17119
rect 22428 17088 22753 17116
rect 22428 17076 22434 17088
rect 22741 17085 22753 17088
rect 22787 17116 22799 17119
rect 22830 17116 22836 17128
rect 22787 17088 22836 17116
rect 22787 17085 22799 17088
rect 22741 17079 22799 17085
rect 22830 17076 22836 17088
rect 22888 17076 22894 17128
rect 20349 17051 20407 17057
rect 20349 17017 20361 17051
rect 20395 17048 20407 17051
rect 20686 17051 20744 17057
rect 20686 17048 20698 17051
rect 20395 17020 20698 17048
rect 20395 17017 20407 17020
rect 20349 17011 20407 17017
rect 20686 17017 20698 17020
rect 20732 17017 20744 17051
rect 20686 17011 20744 17017
rect 22186 17008 22192 17060
rect 22244 17008 22250 17060
rect 22557 17051 22615 17057
rect 22557 17017 22569 17051
rect 22603 17048 22615 17051
rect 22603 17020 22784 17048
rect 22603 17017 22615 17020
rect 22557 17011 22615 17017
rect 22756 16992 22784 17020
rect 21450 16980 21456 16992
rect 19904 16952 21456 16980
rect 21450 16940 21456 16952
rect 21508 16980 21514 16992
rect 21821 16983 21879 16989
rect 21821 16980 21833 16983
rect 21508 16952 21833 16980
rect 21508 16940 21514 16952
rect 21821 16949 21833 16952
rect 21867 16949 21879 16983
rect 21821 16943 21879 16949
rect 22738 16940 22744 16992
rect 22796 16940 22802 16992
rect 552 16890 23368 16912
rect 552 16838 4322 16890
rect 4374 16838 4386 16890
rect 4438 16838 4450 16890
rect 4502 16838 4514 16890
rect 4566 16838 4578 16890
rect 4630 16838 23368 16890
rect 552 16816 23368 16838
rect 3697 16779 3755 16785
rect 3697 16745 3709 16779
rect 3743 16776 3755 16779
rect 4154 16776 4160 16788
rect 3743 16748 4160 16776
rect 3743 16745 3755 16748
rect 3697 16739 3755 16745
rect 4154 16736 4160 16748
rect 4212 16736 4218 16788
rect 4249 16779 4307 16785
rect 4249 16745 4261 16779
rect 4295 16776 4307 16779
rect 5442 16776 5448 16788
rect 4295 16748 5448 16776
rect 4295 16745 4307 16748
rect 4249 16739 4307 16745
rect 5442 16736 5448 16748
rect 5500 16736 5506 16788
rect 7653 16779 7711 16785
rect 7653 16745 7665 16779
rect 7699 16776 7711 16779
rect 9674 16776 9680 16788
rect 7699 16748 9680 16776
rect 7699 16745 7711 16748
rect 7653 16739 7711 16745
rect 9674 16736 9680 16748
rect 9732 16736 9738 16788
rect 11514 16736 11520 16788
rect 11572 16736 11578 16788
rect 12342 16736 12348 16788
rect 12400 16776 12406 16788
rect 15378 16776 15384 16788
rect 12400 16748 15384 16776
rect 12400 16736 12406 16748
rect 15378 16736 15384 16748
rect 15436 16736 15442 16788
rect 16850 16776 16856 16788
rect 15948 16748 16856 16776
rect 2961 16711 3019 16717
rect 2961 16677 2973 16711
rect 3007 16708 3019 16711
rect 3007 16680 3556 16708
rect 3007 16677 3019 16680
rect 2961 16671 3019 16677
rect 3528 16652 3556 16680
rect 3896 16680 4568 16708
rect 3896 16652 3924 16680
rect 2866 16600 2872 16652
rect 2924 16600 2930 16652
rect 3142 16600 3148 16652
rect 3200 16600 3206 16652
rect 3329 16643 3387 16649
rect 3329 16609 3341 16643
rect 3375 16609 3387 16643
rect 3329 16603 3387 16609
rect 3421 16643 3479 16649
rect 3421 16609 3433 16643
rect 3467 16609 3479 16643
rect 3421 16603 3479 16609
rect 3050 16532 3056 16584
rect 3108 16572 3114 16584
rect 3344 16572 3372 16603
rect 3108 16544 3372 16572
rect 3436 16572 3464 16603
rect 3510 16600 3516 16652
rect 3568 16600 3574 16652
rect 3789 16643 3847 16649
rect 3789 16609 3801 16643
rect 3835 16640 3847 16643
rect 3878 16640 3884 16652
rect 3835 16612 3884 16640
rect 3835 16609 3847 16612
rect 3789 16603 3847 16609
rect 3878 16600 3884 16612
rect 3936 16600 3942 16652
rect 3973 16643 4031 16649
rect 3973 16609 3985 16643
rect 4019 16609 4031 16643
rect 3973 16603 4031 16609
rect 3988 16572 4016 16603
rect 4062 16600 4068 16652
rect 4120 16640 4126 16652
rect 4540 16649 4568 16680
rect 7006 16668 7012 16720
rect 7064 16708 7070 16720
rect 7285 16711 7343 16717
rect 7285 16708 7297 16711
rect 7064 16680 7297 16708
rect 7064 16668 7070 16680
rect 7285 16677 7297 16680
rect 7331 16677 7343 16711
rect 7285 16671 7343 16677
rect 7742 16668 7748 16720
rect 7800 16708 7806 16720
rect 8110 16708 8116 16720
rect 7800 16680 8116 16708
rect 7800 16668 7806 16680
rect 8110 16668 8116 16680
rect 8168 16708 8174 16720
rect 8205 16711 8263 16717
rect 8205 16708 8217 16711
rect 8168 16680 8217 16708
rect 8168 16668 8174 16680
rect 8205 16677 8217 16680
rect 8251 16677 8263 16711
rect 8205 16671 8263 16677
rect 8294 16668 8300 16720
rect 8352 16708 8358 16720
rect 8405 16711 8463 16717
rect 8405 16708 8417 16711
rect 8352 16680 8417 16708
rect 8352 16668 8358 16680
rect 8405 16677 8417 16680
rect 8451 16677 8463 16711
rect 11054 16708 11060 16720
rect 8405 16671 8463 16677
rect 10428 16680 11060 16708
rect 4341 16643 4399 16649
rect 4341 16640 4353 16643
rect 4120 16612 4353 16640
rect 4120 16600 4126 16612
rect 4341 16609 4353 16612
rect 4387 16609 4399 16643
rect 4341 16603 4399 16609
rect 4525 16643 4583 16649
rect 4525 16609 4537 16643
rect 4571 16609 4583 16643
rect 4525 16603 4583 16609
rect 4893 16643 4951 16649
rect 4893 16609 4905 16643
rect 4939 16640 4951 16643
rect 5258 16640 5264 16652
rect 4939 16612 5264 16640
rect 4939 16609 4951 16612
rect 4893 16603 4951 16609
rect 4614 16572 4620 16584
rect 3436 16544 3556 16572
rect 3988 16544 4620 16572
rect 3108 16532 3114 16544
rect 3528 16516 3556 16544
rect 4614 16532 4620 16544
rect 4672 16572 4678 16584
rect 4908 16572 4936 16603
rect 5258 16600 5264 16612
rect 5316 16600 5322 16652
rect 5537 16643 5595 16649
rect 5537 16609 5549 16643
rect 5583 16640 5595 16643
rect 6270 16640 6276 16652
rect 5583 16612 6276 16640
rect 5583 16609 5595 16612
rect 5537 16603 5595 16609
rect 6270 16600 6276 16612
rect 6328 16600 6334 16652
rect 7098 16600 7104 16652
rect 7156 16640 7162 16652
rect 7193 16643 7251 16649
rect 7193 16640 7205 16643
rect 7156 16612 7205 16640
rect 7156 16600 7162 16612
rect 7193 16609 7205 16612
rect 7239 16609 7251 16643
rect 7193 16603 7251 16609
rect 7466 16600 7472 16652
rect 7524 16600 7530 16652
rect 10428 16649 10456 16680
rect 11054 16668 11060 16680
rect 11112 16708 11118 16720
rect 12621 16711 12679 16717
rect 12621 16708 12633 16711
rect 11112 16680 11560 16708
rect 11112 16668 11118 16680
rect 11532 16649 11560 16680
rect 11992 16680 12633 16708
rect 11992 16649 12020 16680
rect 12621 16677 12633 16680
rect 12667 16677 12679 16711
rect 12621 16671 12679 16677
rect 12805 16711 12863 16717
rect 12805 16677 12817 16711
rect 12851 16708 12863 16711
rect 13630 16708 13636 16720
rect 12851 16680 13636 16708
rect 12851 16677 12863 16680
rect 12805 16671 12863 16677
rect 13630 16668 13636 16680
rect 13688 16668 13694 16720
rect 13998 16668 14004 16720
rect 14056 16668 14062 16720
rect 15194 16708 15200 16720
rect 15028 16680 15200 16708
rect 10413 16643 10471 16649
rect 10413 16609 10425 16643
rect 10459 16609 10471 16643
rect 11379 16643 11437 16649
rect 11379 16640 11391 16643
rect 10413 16603 10471 16609
rect 10520 16612 11391 16640
rect 4672 16544 4936 16572
rect 4672 16532 4678 16544
rect 6454 16532 6460 16584
rect 6512 16532 6518 16584
rect 7009 16575 7067 16581
rect 7009 16541 7021 16575
rect 7055 16541 7067 16575
rect 7009 16535 7067 16541
rect 3510 16464 3516 16516
rect 3568 16464 3574 16516
rect 7024 16504 7052 16535
rect 9674 16532 9680 16584
rect 9732 16572 9738 16584
rect 10520 16581 10548 16612
rect 11379 16609 11391 16612
rect 11425 16609 11437 16643
rect 11379 16603 11437 16609
rect 11517 16643 11575 16649
rect 11517 16609 11529 16643
rect 11563 16609 11575 16643
rect 11517 16603 11575 16609
rect 11977 16643 12035 16649
rect 11977 16609 11989 16643
rect 12023 16609 12035 16643
rect 12158 16640 12164 16652
rect 11977 16603 12035 16609
rect 12084 16612 12164 16640
rect 10505 16575 10563 16581
rect 10505 16572 10517 16575
rect 9732 16544 10517 16572
rect 9732 16532 9738 16544
rect 10505 16541 10517 16544
rect 10551 16541 10563 16575
rect 10505 16535 10563 16541
rect 10962 16532 10968 16584
rect 11020 16532 11026 16584
rect 7742 16504 7748 16516
rect 7024 16476 7748 16504
rect 7742 16464 7748 16476
rect 7800 16504 7806 16516
rect 8846 16504 8852 16516
rect 7800 16476 8852 16504
rect 7800 16464 7806 16476
rect 8846 16464 8852 16476
rect 8904 16464 8910 16516
rect 10781 16507 10839 16513
rect 10781 16473 10793 16507
rect 10827 16504 10839 16507
rect 11992 16504 12020 16603
rect 12084 16581 12112 16612
rect 12158 16600 12164 16612
rect 12216 16640 12222 16652
rect 12437 16643 12495 16649
rect 12437 16640 12449 16643
rect 12216 16612 12449 16640
rect 12216 16600 12222 16612
rect 12437 16609 12449 16612
rect 12483 16609 12495 16643
rect 12437 16603 12495 16609
rect 13722 16600 13728 16652
rect 13780 16600 13786 16652
rect 13817 16643 13875 16649
rect 13817 16609 13829 16643
rect 13863 16640 13875 16643
rect 13906 16640 13912 16652
rect 13863 16612 13912 16640
rect 13863 16609 13875 16612
rect 13817 16603 13875 16609
rect 13906 16600 13912 16612
rect 13964 16600 13970 16652
rect 15028 16640 15056 16680
rect 15194 16668 15200 16680
rect 15252 16668 15258 16720
rect 14108 16612 15056 16640
rect 12069 16575 12127 16581
rect 12069 16541 12081 16575
rect 12115 16541 12127 16575
rect 12069 16535 12127 16541
rect 12342 16532 12348 16584
rect 12400 16532 12406 16584
rect 14108 16572 14136 16612
rect 15102 16600 15108 16652
rect 15160 16640 15166 16652
rect 15289 16643 15347 16649
rect 15160 16612 15240 16640
rect 15160 16600 15166 16612
rect 14016 16544 14136 16572
rect 15212 16572 15240 16612
rect 15289 16609 15301 16643
rect 15335 16640 15347 16643
rect 15565 16643 15623 16649
rect 15565 16640 15577 16643
rect 15335 16612 15577 16640
rect 15335 16609 15347 16612
rect 15289 16603 15347 16609
rect 15565 16609 15577 16612
rect 15611 16640 15623 16643
rect 15654 16640 15660 16652
rect 15611 16612 15660 16640
rect 15611 16609 15623 16612
rect 15565 16603 15623 16609
rect 15654 16600 15660 16612
rect 15712 16600 15718 16652
rect 15948 16640 15976 16748
rect 16850 16736 16856 16748
rect 16908 16736 16914 16788
rect 18138 16736 18144 16788
rect 18196 16736 18202 16788
rect 18414 16736 18420 16788
rect 18472 16736 18478 16788
rect 18601 16779 18659 16785
rect 18601 16745 18613 16779
rect 18647 16776 18659 16779
rect 18966 16776 18972 16788
rect 18647 16748 18972 16776
rect 18647 16745 18659 16748
rect 18601 16739 18659 16745
rect 18966 16736 18972 16748
rect 19024 16736 19030 16788
rect 19150 16736 19156 16788
rect 19208 16776 19214 16788
rect 20073 16779 20131 16785
rect 20073 16776 20085 16779
rect 19208 16748 20085 16776
rect 19208 16736 19214 16748
rect 20073 16745 20085 16748
rect 20119 16745 20131 16779
rect 20073 16739 20131 16745
rect 22830 16736 22836 16788
rect 22888 16736 22894 16788
rect 16022 16668 16028 16720
rect 16080 16708 16086 16720
rect 18432 16708 18460 16736
rect 18874 16708 18880 16720
rect 16080 16680 16620 16708
rect 16080 16668 16086 16680
rect 16592 16649 16620 16680
rect 17788 16680 18460 16708
rect 18708 16680 18880 16708
rect 16117 16643 16175 16649
rect 16117 16640 16129 16643
rect 15948 16612 16129 16640
rect 16117 16609 16129 16612
rect 16163 16609 16175 16643
rect 16117 16603 16175 16609
rect 16301 16643 16359 16649
rect 16301 16609 16313 16643
rect 16347 16609 16359 16643
rect 16301 16603 16359 16609
rect 16577 16643 16635 16649
rect 16577 16609 16589 16643
rect 16623 16609 16635 16643
rect 16577 16603 16635 16609
rect 15473 16575 15531 16581
rect 15473 16572 15485 16575
rect 15212 16544 15485 16572
rect 14016 16513 14044 16544
rect 15473 16541 15485 16544
rect 15519 16541 15531 16575
rect 15473 16535 15531 16541
rect 15838 16532 15844 16584
rect 15896 16572 15902 16584
rect 16316 16572 16344 16603
rect 17126 16600 17132 16652
rect 17184 16600 17190 16652
rect 17310 16600 17316 16652
rect 17368 16600 17374 16652
rect 17788 16649 17816 16680
rect 17497 16643 17555 16649
rect 17497 16609 17509 16643
rect 17543 16609 17555 16643
rect 17497 16603 17555 16609
rect 17773 16643 17831 16649
rect 17773 16609 17785 16643
rect 17819 16609 17831 16643
rect 17773 16603 17831 16609
rect 15896 16544 16344 16572
rect 16761 16575 16819 16581
rect 15896 16532 15902 16544
rect 16761 16541 16773 16575
rect 16807 16572 16819 16575
rect 16942 16572 16948 16584
rect 16807 16544 16948 16572
rect 16807 16541 16819 16544
rect 16761 16535 16819 16541
rect 16942 16532 16948 16544
rect 17000 16572 17006 16584
rect 17512 16572 17540 16603
rect 17862 16600 17868 16652
rect 17920 16640 17926 16652
rect 18049 16643 18107 16649
rect 18049 16640 18061 16643
rect 17920 16612 18061 16640
rect 17920 16600 17926 16612
rect 18049 16609 18061 16612
rect 18095 16640 18107 16643
rect 18233 16643 18291 16649
rect 18233 16640 18245 16643
rect 18095 16612 18245 16640
rect 18095 16609 18107 16612
rect 18049 16603 18107 16609
rect 18233 16609 18245 16612
rect 18279 16609 18291 16643
rect 18233 16603 18291 16609
rect 18322 16600 18328 16652
rect 18380 16640 18386 16652
rect 18417 16643 18475 16649
rect 18417 16640 18429 16643
rect 18380 16612 18429 16640
rect 18380 16600 18386 16612
rect 18417 16609 18429 16612
rect 18463 16609 18475 16643
rect 18417 16603 18475 16609
rect 18708 16581 18736 16680
rect 18874 16668 18880 16680
rect 18932 16708 18938 16720
rect 20438 16708 20444 16720
rect 18932 16680 20444 16708
rect 18932 16668 18938 16680
rect 20438 16668 20444 16680
rect 20496 16668 20502 16720
rect 22646 16708 22652 16720
rect 21468 16680 22652 16708
rect 18960 16643 19018 16649
rect 18960 16609 18972 16643
rect 19006 16640 19018 16643
rect 19242 16640 19248 16652
rect 19006 16612 19248 16640
rect 19006 16609 19018 16612
rect 18960 16603 19018 16609
rect 19242 16600 19248 16612
rect 19300 16600 19306 16652
rect 21174 16600 21180 16652
rect 21232 16640 21238 16652
rect 21468 16649 21496 16680
rect 22646 16668 22652 16680
rect 22704 16668 22710 16720
rect 21726 16649 21732 16652
rect 21453 16643 21511 16649
rect 21453 16640 21465 16643
rect 21232 16612 21465 16640
rect 21232 16600 21238 16612
rect 21453 16609 21465 16612
rect 21499 16609 21511 16643
rect 21720 16640 21732 16649
rect 21687 16612 21732 16640
rect 21453 16603 21511 16609
rect 21720 16603 21732 16612
rect 21726 16600 21732 16603
rect 21784 16600 21790 16652
rect 18693 16575 18751 16581
rect 18693 16572 18705 16575
rect 17000 16544 17540 16572
rect 18248 16544 18705 16572
rect 17000 16532 17006 16544
rect 10827 16476 12020 16504
rect 14001 16507 14059 16513
rect 10827 16473 10839 16476
rect 10781 16467 10839 16473
rect 14001 16473 14013 16507
rect 14047 16473 14059 16507
rect 14001 16467 14059 16473
rect 15105 16507 15163 16513
rect 15105 16473 15117 16507
rect 15151 16504 15163 16507
rect 15856 16504 15884 16532
rect 18248 16516 18276 16544
rect 18693 16541 18705 16544
rect 18739 16541 18751 16575
rect 18693 16535 18751 16541
rect 15151 16476 15884 16504
rect 15151 16473 15163 16476
rect 15105 16467 15163 16473
rect 18230 16464 18236 16516
rect 18288 16464 18294 16516
rect 8202 16396 8208 16448
rect 8260 16436 8266 16448
rect 8389 16439 8447 16445
rect 8389 16436 8401 16439
rect 8260 16408 8401 16436
rect 8260 16396 8266 16408
rect 8389 16405 8401 16408
rect 8435 16405 8447 16439
rect 8389 16399 8447 16405
rect 8570 16396 8576 16448
rect 8628 16396 8634 16448
rect 15841 16439 15899 16445
rect 15841 16405 15853 16439
rect 15887 16436 15899 16439
rect 16482 16436 16488 16448
rect 15887 16408 16488 16436
rect 15887 16405 15899 16408
rect 15841 16399 15899 16405
rect 16482 16396 16488 16408
rect 16540 16396 16546 16448
rect 552 16346 23368 16368
rect 552 16294 3662 16346
rect 3714 16294 3726 16346
rect 3778 16294 3790 16346
rect 3842 16294 3854 16346
rect 3906 16294 3918 16346
rect 3970 16294 23368 16346
rect 552 16272 23368 16294
rect 9030 16232 9036 16244
rect 7852 16204 9036 16232
rect 3142 16124 3148 16176
rect 3200 16164 3206 16176
rect 3513 16167 3571 16173
rect 3513 16164 3525 16167
rect 3200 16136 3525 16164
rect 3200 16124 3206 16136
rect 3513 16133 3525 16136
rect 3559 16133 3571 16167
rect 3513 16127 3571 16133
rect 4985 16167 5043 16173
rect 4985 16133 4997 16167
rect 5031 16133 5043 16167
rect 4985 16127 5043 16133
rect 3418 16096 3424 16108
rect 2700 16068 3424 16096
rect 2700 16037 2728 16068
rect 3418 16056 3424 16068
rect 3476 16096 3482 16108
rect 3881 16099 3939 16105
rect 3881 16096 3893 16099
rect 3476 16068 3893 16096
rect 3476 16056 3482 16068
rect 3881 16065 3893 16068
rect 3927 16096 3939 16099
rect 3970 16096 3976 16108
rect 3927 16068 3976 16096
rect 3927 16065 3939 16068
rect 3881 16059 3939 16065
rect 3970 16056 3976 16068
rect 4028 16056 4034 16108
rect 4154 16056 4160 16108
rect 4212 16096 4218 16108
rect 4525 16099 4583 16105
rect 4525 16096 4537 16099
rect 4212 16068 4537 16096
rect 4212 16056 4218 16068
rect 4525 16065 4537 16068
rect 4571 16065 4583 16099
rect 5000 16096 5028 16127
rect 5905 16099 5963 16105
rect 5905 16096 5917 16099
rect 5000 16068 5917 16096
rect 4525 16059 4583 16065
rect 5905 16065 5917 16068
rect 5951 16096 5963 16099
rect 6086 16096 6092 16108
rect 5951 16068 6092 16096
rect 5951 16065 5963 16068
rect 5905 16059 5963 16065
rect 6086 16056 6092 16068
rect 6144 16056 6150 16108
rect 6181 16099 6239 16105
rect 6181 16065 6193 16099
rect 6227 16096 6239 16099
rect 7098 16096 7104 16108
rect 6227 16068 7104 16096
rect 6227 16065 6239 16068
rect 6181 16059 6239 16065
rect 7098 16056 7104 16068
rect 7156 16056 7162 16108
rect 7742 16056 7748 16108
rect 7800 16056 7806 16108
rect 2685 16031 2743 16037
rect 2685 15997 2697 16031
rect 2731 15997 2743 16031
rect 3510 16028 3516 16040
rect 2685 15991 2743 15997
rect 2884 16000 3516 16028
rect 2884 15972 2912 16000
rect 3510 15988 3516 16000
rect 3568 16028 3574 16040
rect 3789 16031 3847 16037
rect 3789 16028 3801 16031
rect 3568 16000 3801 16028
rect 3568 15988 3574 16000
rect 3789 15997 3801 16000
rect 3835 16028 3847 16031
rect 4065 16031 4123 16037
rect 4065 16028 4077 16031
rect 3835 16000 4077 16028
rect 3835 15997 3847 16000
rect 3789 15991 3847 15997
rect 4065 15997 4077 16000
rect 4111 15997 4123 16031
rect 4065 15991 4123 15997
rect 4614 15988 4620 16040
rect 4672 15988 4678 16040
rect 5442 15988 5448 16040
rect 5500 16028 5506 16040
rect 5813 16031 5871 16037
rect 5813 16028 5825 16031
rect 5500 16000 5825 16028
rect 5500 15988 5506 16000
rect 5813 15997 5825 16000
rect 5859 15997 5871 16031
rect 5813 15991 5871 15997
rect 6270 15988 6276 16040
rect 6328 15988 6334 16040
rect 6454 15988 6460 16040
rect 6512 15988 6518 16040
rect 7190 15988 7196 16040
rect 7248 15988 7254 16040
rect 7852 16037 7880 16204
rect 9030 16192 9036 16204
rect 9088 16192 9094 16244
rect 9674 16192 9680 16244
rect 9732 16192 9738 16244
rect 9861 16235 9919 16241
rect 9861 16201 9873 16235
rect 9907 16232 9919 16235
rect 10962 16232 10968 16244
rect 9907 16204 10968 16232
rect 9907 16201 9919 16204
rect 9861 16195 9919 16201
rect 10962 16192 10968 16204
rect 11020 16192 11026 16244
rect 13538 16192 13544 16244
rect 13596 16192 13602 16244
rect 15838 16192 15844 16244
rect 15896 16192 15902 16244
rect 15930 16192 15936 16244
rect 15988 16232 15994 16244
rect 16209 16235 16267 16241
rect 16209 16232 16221 16235
rect 15988 16204 16221 16232
rect 15988 16192 15994 16204
rect 16209 16201 16221 16204
rect 16255 16201 16267 16235
rect 16209 16195 16267 16201
rect 16850 16192 16856 16244
rect 16908 16192 16914 16244
rect 17037 16235 17095 16241
rect 17037 16201 17049 16235
rect 17083 16232 17095 16235
rect 17310 16232 17316 16244
rect 17083 16204 17316 16232
rect 17083 16201 17095 16204
rect 17037 16195 17095 16201
rect 8205 16167 8263 16173
rect 8205 16133 8217 16167
rect 8251 16164 8263 16167
rect 8294 16164 8300 16176
rect 8251 16136 8300 16164
rect 8251 16133 8263 16136
rect 8205 16127 8263 16133
rect 8294 16124 8300 16136
rect 8352 16124 8358 16176
rect 11425 16167 11483 16173
rect 11425 16133 11437 16167
rect 11471 16164 11483 16167
rect 12618 16164 12624 16176
rect 11471 16136 12624 16164
rect 11471 16133 11483 16136
rect 11425 16127 11483 16133
rect 12618 16124 12624 16136
rect 12676 16124 12682 16176
rect 14461 16167 14519 16173
rect 14461 16133 14473 16167
rect 14507 16164 14519 16167
rect 15381 16167 15439 16173
rect 15381 16164 15393 16167
rect 14507 16136 15393 16164
rect 14507 16133 14519 16136
rect 14461 16127 14519 16133
rect 15381 16133 15393 16136
rect 15427 16133 15439 16167
rect 15381 16127 15439 16133
rect 16393 16167 16451 16173
rect 16393 16133 16405 16167
rect 16439 16164 16451 16167
rect 17052 16164 17080 16195
rect 17310 16192 17316 16204
rect 17368 16192 17374 16244
rect 17954 16192 17960 16244
rect 18012 16232 18018 16244
rect 18233 16235 18291 16241
rect 18233 16232 18245 16235
rect 18012 16204 18245 16232
rect 18012 16192 18018 16204
rect 18233 16201 18245 16204
rect 18279 16201 18291 16235
rect 18233 16195 18291 16201
rect 19242 16192 19248 16244
rect 19300 16192 19306 16244
rect 21634 16192 21640 16244
rect 21692 16232 21698 16244
rect 21913 16235 21971 16241
rect 21913 16232 21925 16235
rect 21692 16204 21925 16232
rect 21692 16192 21698 16204
rect 21913 16201 21925 16204
rect 21959 16201 21971 16235
rect 21913 16195 21971 16201
rect 22002 16192 22008 16244
rect 22060 16192 22066 16244
rect 16439 16136 17080 16164
rect 18095 16167 18153 16173
rect 16439 16133 16451 16136
rect 16393 16127 16451 16133
rect 18095 16133 18107 16167
rect 18141 16164 18153 16167
rect 18966 16164 18972 16176
rect 18141 16136 18972 16164
rect 18141 16133 18153 16136
rect 18095 16127 18153 16133
rect 18966 16124 18972 16136
rect 19024 16124 19030 16176
rect 19521 16167 19579 16173
rect 19521 16164 19533 16167
rect 19076 16136 19533 16164
rect 8018 16056 8024 16108
rect 8076 16096 8082 16108
rect 9217 16099 9275 16105
rect 9217 16096 9229 16099
rect 8076 16068 9229 16096
rect 8076 16056 8082 16068
rect 9217 16065 9229 16068
rect 9263 16096 9275 16099
rect 9263 16068 9812 16096
rect 9263 16065 9275 16068
rect 9217 16059 9275 16065
rect 7837 16031 7895 16037
rect 7837 15997 7849 16031
rect 7883 15997 7895 16031
rect 7837 15991 7895 15997
rect 8573 16031 8631 16037
rect 8573 15997 8585 16031
rect 8619 16028 8631 16031
rect 8662 16028 8668 16040
rect 8619 16000 8668 16028
rect 8619 15997 8631 16000
rect 8573 15991 8631 15997
rect 8662 15988 8668 16000
rect 8720 15988 8726 16040
rect 8846 15988 8852 16040
rect 8904 15988 8910 16040
rect 9030 15988 9036 16040
rect 9088 15988 9094 16040
rect 9784 16037 9812 16068
rect 13998 16056 14004 16108
rect 14056 16096 14062 16108
rect 14553 16099 14611 16105
rect 14553 16096 14565 16099
rect 14056 16068 14565 16096
rect 14056 16056 14062 16068
rect 14553 16065 14565 16068
rect 14599 16065 14611 16099
rect 14553 16059 14611 16065
rect 15657 16099 15715 16105
rect 15657 16065 15669 16099
rect 15703 16096 15715 16099
rect 16022 16096 16028 16108
rect 15703 16068 16028 16096
rect 15703 16065 15715 16068
rect 15657 16059 15715 16065
rect 16022 16056 16028 16068
rect 16080 16056 16086 16108
rect 19076 16096 19104 16136
rect 19521 16133 19533 16136
rect 19567 16164 19579 16167
rect 19886 16164 19892 16176
rect 19567 16136 19892 16164
rect 19567 16133 19579 16136
rect 19521 16127 19579 16133
rect 19886 16124 19892 16136
rect 19944 16124 19950 16176
rect 22278 16164 22284 16176
rect 21744 16136 22284 16164
rect 21744 16105 21772 16136
rect 22278 16124 22284 16136
rect 22336 16124 22342 16176
rect 17972 16068 19104 16096
rect 17972 16040 18000 16068
rect 9309 16031 9367 16037
rect 9309 15997 9321 16031
rect 9355 15997 9367 16031
rect 9309 15991 9367 15997
rect 9769 16031 9827 16037
rect 9769 15997 9781 16031
rect 9815 15997 9827 16031
rect 9769 15991 9827 15997
rect 9953 16031 10011 16037
rect 9953 15997 9965 16031
rect 9999 15997 10011 16031
rect 9953 15991 10011 15997
rect 2866 15920 2872 15972
rect 2924 15920 2930 15972
rect 2958 15920 2964 15972
rect 3016 15960 3022 15972
rect 3237 15963 3295 15969
rect 3237 15960 3249 15963
rect 3016 15932 3249 15960
rect 3016 15920 3022 15932
rect 3237 15929 3249 15932
rect 3283 15960 3295 15963
rect 3602 15960 3608 15972
rect 3283 15932 3608 15960
rect 3283 15929 3295 15932
rect 3237 15923 3295 15929
rect 3602 15920 3608 15932
rect 3660 15920 3666 15972
rect 3694 15920 3700 15972
rect 3752 15960 3758 15972
rect 4632 15960 4660 15988
rect 9324 15960 9352 15991
rect 9968 15960 9996 15991
rect 10962 15988 10968 16040
rect 11020 16028 11026 16040
rect 11149 16031 11207 16037
rect 11149 16028 11161 16031
rect 11020 16000 11161 16028
rect 11020 15988 11026 16000
rect 11149 15997 11161 16000
rect 11195 15997 11207 16031
rect 11149 15991 11207 15997
rect 12802 15988 12808 16040
rect 12860 16028 12866 16040
rect 13173 16031 13231 16037
rect 13173 16028 13185 16031
rect 12860 16000 13185 16028
rect 12860 15988 12866 16000
rect 13173 15997 13185 16000
rect 13219 16028 13231 16031
rect 13262 16028 13268 16040
rect 13219 16000 13268 16028
rect 13219 15997 13231 16000
rect 13173 15991 13231 15997
rect 13262 15988 13268 16000
rect 13320 15988 13326 16040
rect 13357 16031 13415 16037
rect 13357 15997 13369 16031
rect 13403 16028 13415 16031
rect 13446 16028 13452 16040
rect 13403 16000 13452 16028
rect 13403 15997 13415 16000
rect 13357 15991 13415 15997
rect 13446 15988 13452 16000
rect 13504 15988 13510 16040
rect 13722 15988 13728 16040
rect 13780 15988 13786 16040
rect 13906 15988 13912 16040
rect 13964 15988 13970 16040
rect 15378 15988 15384 16040
rect 15436 16028 15442 16040
rect 15933 16031 15991 16037
rect 15933 16028 15945 16031
rect 15436 16000 15945 16028
rect 15436 15988 15442 16000
rect 15933 15997 15945 16000
rect 15979 15997 15991 16031
rect 15933 15991 15991 15997
rect 3752 15932 4660 15960
rect 7576 15932 9996 15960
rect 3752 15920 3758 15932
rect 3050 15852 3056 15904
rect 3108 15852 3114 15904
rect 3786 15852 3792 15904
rect 3844 15892 3850 15904
rect 4157 15895 4215 15901
rect 4157 15892 4169 15895
rect 3844 15864 4169 15892
rect 3844 15852 3850 15864
rect 4157 15861 4169 15864
rect 4203 15861 4215 15895
rect 4157 15855 4215 15861
rect 6362 15852 6368 15904
rect 6420 15852 6426 15904
rect 7576 15901 7604 15932
rect 11054 15920 11060 15972
rect 11112 15960 11118 15972
rect 11241 15963 11299 15969
rect 11241 15960 11253 15963
rect 11112 15932 11253 15960
rect 11112 15920 11118 15932
rect 11241 15929 11253 15932
rect 11287 15929 11299 15963
rect 11241 15923 11299 15929
rect 11425 15963 11483 15969
rect 11425 15929 11437 15963
rect 11471 15960 11483 15963
rect 11606 15960 11612 15972
rect 11471 15932 11612 15960
rect 11471 15929 11483 15932
rect 11425 15923 11483 15929
rect 11606 15920 11612 15932
rect 11664 15920 11670 15972
rect 14185 15963 14243 15969
rect 14185 15960 14197 15963
rect 13188 15932 14197 15960
rect 13188 15904 13216 15932
rect 14185 15929 14197 15932
rect 14231 15929 14243 15963
rect 14185 15923 14243 15929
rect 14645 15963 14703 15969
rect 14645 15929 14657 15963
rect 14691 15929 14703 15963
rect 15948 15960 15976 15991
rect 16482 15988 16488 16040
rect 16540 15988 16546 16040
rect 16758 15988 16764 16040
rect 16816 15988 16822 16040
rect 16942 15988 16948 16040
rect 17000 16028 17006 16040
rect 17037 16031 17095 16037
rect 17037 16028 17049 16031
rect 17000 16000 17049 16028
rect 17000 15988 17006 16000
rect 17037 15997 17049 16000
rect 17083 15997 17095 16031
rect 17037 15991 17095 15997
rect 17126 15988 17132 16040
rect 17184 15988 17190 16040
rect 17954 15988 17960 16040
rect 18012 15988 18018 16040
rect 18414 15988 18420 16040
rect 18472 15988 18478 16040
rect 18690 15988 18696 16040
rect 18748 15988 18754 16040
rect 18782 15988 18788 16040
rect 18840 16028 18846 16040
rect 19076 16037 19104 16068
rect 21729 16099 21787 16105
rect 21729 16065 21741 16099
rect 21775 16065 21787 16099
rect 21729 16059 21787 16065
rect 21821 16099 21879 16105
rect 21821 16065 21833 16099
rect 21867 16096 21879 16099
rect 22186 16096 22192 16108
rect 21867 16068 22192 16096
rect 21867 16065 21879 16068
rect 21821 16059 21879 16065
rect 18877 16031 18935 16037
rect 18877 16028 18889 16031
rect 18840 16000 18889 16028
rect 18840 15988 18846 16000
rect 18877 15997 18889 16000
rect 18923 15997 18935 16031
rect 18877 15991 18935 15997
rect 19061 16031 19119 16037
rect 19061 15997 19073 16031
rect 19107 15997 19119 16031
rect 19061 15991 19119 15997
rect 19337 16031 19395 16037
rect 19337 15997 19349 16031
rect 19383 16028 19395 16031
rect 19518 16028 19524 16040
rect 19383 16000 19524 16028
rect 19383 15997 19395 16000
rect 19337 15991 19395 15997
rect 19518 15988 19524 16000
rect 19576 15988 19582 16040
rect 21450 15988 21456 16040
rect 21508 15988 21514 16040
rect 21542 15988 21548 16040
rect 21600 15988 21606 16040
rect 16025 15963 16083 15969
rect 16025 15960 16037 15963
rect 15948 15932 16037 15960
rect 14645 15923 14703 15929
rect 16025 15929 16037 15932
rect 16071 15929 16083 15963
rect 16025 15923 16083 15929
rect 16241 15963 16299 15969
rect 16241 15929 16253 15963
rect 16287 15960 16299 15963
rect 16574 15960 16580 15972
rect 16287 15932 16580 15960
rect 16287 15929 16299 15932
rect 16241 15923 16299 15929
rect 7561 15895 7619 15901
rect 7561 15861 7573 15895
rect 7607 15861 7619 15895
rect 7561 15855 7619 15861
rect 8386 15852 8392 15904
rect 8444 15852 8450 15904
rect 13170 15852 13176 15904
rect 13228 15852 13234 15904
rect 13265 15895 13323 15901
rect 13265 15861 13277 15895
rect 13311 15892 13323 15895
rect 13446 15892 13452 15904
rect 13311 15864 13452 15892
rect 13311 15861 13323 15864
rect 13265 15855 13323 15861
rect 13446 15852 13452 15864
rect 13504 15852 13510 15904
rect 13722 15852 13728 15904
rect 13780 15892 13786 15904
rect 14277 15895 14335 15901
rect 14277 15892 14289 15895
rect 13780 15864 14289 15892
rect 13780 15852 13786 15864
rect 14277 15861 14289 15864
rect 14323 15861 14335 15895
rect 14660 15892 14688 15923
rect 16574 15920 16580 15932
rect 16632 15920 16638 15972
rect 17144 15892 17172 15988
rect 18969 15963 19027 15969
rect 18969 15929 18981 15963
rect 19015 15960 19027 15963
rect 19150 15960 19156 15972
rect 19015 15932 19156 15960
rect 19015 15929 19027 15932
rect 18969 15923 19027 15929
rect 19150 15920 19156 15932
rect 19208 15920 19214 15972
rect 19536 15960 19564 15988
rect 21836 15960 21864 16059
rect 22186 16056 22192 16068
rect 22244 16056 22250 16108
rect 22094 15988 22100 16040
rect 22152 15988 22158 16040
rect 19536 15932 21864 15960
rect 14660 15864 17172 15892
rect 17405 15895 17463 15901
rect 14277 15855 14335 15861
rect 17405 15861 17417 15895
rect 17451 15892 17463 15895
rect 18322 15892 18328 15904
rect 17451 15864 18328 15892
rect 17451 15861 17463 15864
rect 17405 15855 17463 15861
rect 18322 15852 18328 15864
rect 18380 15852 18386 15904
rect 18417 15895 18475 15901
rect 18417 15861 18429 15895
rect 18463 15892 18475 15895
rect 18506 15892 18512 15904
rect 18463 15864 18512 15892
rect 18463 15861 18475 15864
rect 18417 15855 18475 15861
rect 18506 15852 18512 15864
rect 18564 15852 18570 15904
rect 21726 15852 21732 15904
rect 21784 15852 21790 15904
rect 552 15802 23368 15824
rect 552 15750 4322 15802
rect 4374 15750 4386 15802
rect 4438 15750 4450 15802
rect 4502 15750 4514 15802
rect 4566 15750 4578 15802
rect 4630 15750 23368 15802
rect 552 15728 23368 15750
rect 3050 15648 3056 15700
rect 3108 15688 3114 15700
rect 3329 15691 3387 15697
rect 3329 15688 3341 15691
rect 3108 15660 3341 15688
rect 3108 15648 3114 15660
rect 3329 15657 3341 15660
rect 3375 15688 3387 15691
rect 3375 15660 4292 15688
rect 3375 15657 3387 15660
rect 3329 15651 3387 15657
rect 3694 15629 3700 15632
rect 3671 15623 3700 15629
rect 3671 15589 3683 15623
rect 3671 15583 3700 15589
rect 3694 15580 3700 15583
rect 3752 15580 3758 15632
rect 3786 15580 3792 15632
rect 3844 15580 3850 15632
rect 4264 15629 4292 15660
rect 8018 15648 8024 15700
rect 8076 15648 8082 15700
rect 8294 15648 8300 15700
rect 8352 15648 8358 15700
rect 11606 15648 11612 15700
rect 11664 15648 11670 15700
rect 13541 15691 13599 15697
rect 13541 15657 13553 15691
rect 13587 15688 13599 15691
rect 13722 15688 13728 15700
rect 13587 15660 13728 15688
rect 13587 15657 13599 15660
rect 13541 15651 13599 15657
rect 13722 15648 13728 15660
rect 13780 15648 13786 15700
rect 21818 15648 21824 15700
rect 21876 15688 21882 15700
rect 22557 15691 22615 15697
rect 22557 15688 22569 15691
rect 21876 15660 22569 15688
rect 21876 15648 21882 15660
rect 22557 15657 22569 15660
rect 22603 15657 22615 15691
rect 22557 15651 22615 15657
rect 4249 15623 4307 15629
rect 4249 15589 4261 15623
rect 4295 15589 4307 15623
rect 4249 15583 4307 15589
rect 4341 15623 4399 15629
rect 4341 15589 4353 15623
rect 4387 15620 4399 15623
rect 6454 15620 6460 15632
rect 4387 15592 6460 15620
rect 4387 15589 4399 15592
rect 4341 15583 4399 15589
rect 6454 15580 6460 15592
rect 6512 15580 6518 15632
rect 7190 15580 7196 15632
rect 7248 15620 7254 15632
rect 8312 15620 8340 15648
rect 8573 15623 8631 15629
rect 8573 15620 8585 15623
rect 7248 15592 7972 15620
rect 8312 15592 8585 15620
rect 7248 15580 7254 15592
rect 3142 15512 3148 15564
rect 3200 15552 3206 15564
rect 3421 15555 3479 15561
rect 3421 15552 3433 15555
rect 3200 15524 3433 15552
rect 3200 15512 3206 15524
rect 3421 15521 3433 15524
rect 3467 15552 3479 15555
rect 3467 15524 3648 15552
rect 3467 15521 3479 15524
rect 3421 15515 3479 15521
rect 2958 15444 2964 15496
rect 3016 15444 3022 15496
rect 3513 15487 3571 15493
rect 3513 15453 3525 15487
rect 3559 15453 3571 15487
rect 3620 15484 3648 15524
rect 3878 15512 3884 15564
rect 3936 15512 3942 15564
rect 3970 15512 3976 15564
rect 4028 15512 4034 15564
rect 4617 15555 4675 15561
rect 4617 15552 4629 15555
rect 4080 15524 4629 15552
rect 4080 15484 4108 15524
rect 4617 15521 4629 15524
rect 4663 15521 4675 15555
rect 4617 15515 4675 15521
rect 4706 15512 4712 15564
rect 4764 15552 4770 15564
rect 4801 15555 4859 15561
rect 4801 15552 4813 15555
rect 4764 15524 4813 15552
rect 4764 15512 4770 15524
rect 4801 15521 4813 15524
rect 4847 15521 4859 15555
rect 4801 15515 4859 15521
rect 7742 15512 7748 15564
rect 7800 15512 7806 15564
rect 7944 15561 7972 15592
rect 8573 15589 8585 15592
rect 8619 15589 8631 15623
rect 8573 15583 8631 15589
rect 11348 15592 11928 15620
rect 11348 15564 11376 15592
rect 7929 15555 7987 15561
rect 7929 15521 7941 15555
rect 7975 15521 7987 15555
rect 7929 15515 7987 15521
rect 8202 15512 8208 15564
rect 8260 15552 8266 15564
rect 8297 15555 8355 15561
rect 8297 15552 8309 15555
rect 8260 15524 8309 15552
rect 8260 15512 8266 15524
rect 8297 15521 8309 15524
rect 8343 15521 8355 15555
rect 8297 15515 8355 15521
rect 8389 15555 8447 15561
rect 8389 15521 8401 15555
rect 8435 15521 8447 15555
rect 8389 15515 8447 15521
rect 3620 15456 4108 15484
rect 3513 15447 3571 15453
rect 3145 15419 3203 15425
rect 3145 15385 3157 15419
rect 3191 15416 3203 15419
rect 3528 15416 3556 15447
rect 8110 15444 8116 15496
rect 8168 15484 8174 15496
rect 8404 15484 8432 15515
rect 11330 15512 11336 15564
rect 11388 15512 11394 15564
rect 11900 15561 11928 15592
rect 13280 15592 14136 15620
rect 13280 15564 13308 15592
rect 11793 15555 11851 15561
rect 11793 15521 11805 15555
rect 11839 15521 11851 15555
rect 11793 15515 11851 15521
rect 11885 15555 11943 15561
rect 11885 15521 11897 15555
rect 11931 15521 11943 15555
rect 11885 15515 11943 15521
rect 8168 15456 8432 15484
rect 8168 15444 8174 15456
rect 10962 15444 10968 15496
rect 11020 15444 11026 15496
rect 11238 15444 11244 15496
rect 11296 15484 11302 15496
rect 11808 15484 11836 15515
rect 13262 15512 13268 15564
rect 13320 15512 13326 15564
rect 13446 15512 13452 15564
rect 13504 15552 13510 15564
rect 13725 15555 13783 15561
rect 13725 15552 13737 15555
rect 13504 15524 13737 15552
rect 13504 15512 13510 15524
rect 13725 15521 13737 15524
rect 13771 15521 13783 15555
rect 13725 15515 13783 15521
rect 13814 15512 13820 15564
rect 13872 15552 13878 15564
rect 14108 15561 14136 15592
rect 15396 15592 15884 15620
rect 15396 15564 15424 15592
rect 13909 15555 13967 15561
rect 13909 15552 13921 15555
rect 13872 15524 13921 15552
rect 13872 15512 13878 15524
rect 13909 15521 13921 15524
rect 13955 15521 13967 15555
rect 13909 15515 13967 15521
rect 14001 15555 14059 15561
rect 14001 15521 14013 15555
rect 14047 15521 14059 15555
rect 14001 15515 14059 15521
rect 14093 15555 14151 15561
rect 14093 15521 14105 15555
rect 14139 15521 14151 15555
rect 14093 15515 14151 15521
rect 14277 15555 14335 15561
rect 14277 15521 14289 15555
rect 14323 15521 14335 15555
rect 14277 15515 14335 15521
rect 11296 15456 11836 15484
rect 11296 15444 11302 15456
rect 13354 15444 13360 15496
rect 13412 15444 13418 15496
rect 14016 15484 14044 15515
rect 14185 15487 14243 15493
rect 14185 15484 14197 15487
rect 14016 15456 14197 15484
rect 14185 15453 14197 15456
rect 14231 15453 14243 15487
rect 14185 15447 14243 15453
rect 4706 15416 4712 15428
rect 3191 15388 4712 15416
rect 3191 15385 3203 15388
rect 3145 15379 3203 15385
rect 4706 15376 4712 15388
rect 4764 15376 4770 15428
rect 6362 15376 6368 15428
rect 6420 15416 6426 15428
rect 8205 15419 8263 15425
rect 8205 15416 8217 15419
rect 6420 15388 8217 15416
rect 6420 15376 6426 15388
rect 8205 15385 8217 15388
rect 8251 15416 8263 15419
rect 8662 15416 8668 15428
rect 8251 15388 8668 15416
rect 8251 15385 8263 15388
rect 8205 15379 8263 15385
rect 8662 15376 8668 15388
rect 8720 15376 8726 15428
rect 12894 15376 12900 15428
rect 12952 15376 12958 15428
rect 13372 15416 13400 15444
rect 14292 15416 14320 15515
rect 15010 15512 15016 15564
rect 15068 15512 15074 15564
rect 15194 15512 15200 15564
rect 15252 15512 15258 15564
rect 15289 15555 15347 15561
rect 15289 15521 15301 15555
rect 15335 15552 15347 15555
rect 15378 15552 15384 15564
rect 15335 15524 15384 15552
rect 15335 15521 15347 15524
rect 15289 15515 15347 15521
rect 15378 15512 15384 15524
rect 15436 15512 15442 15564
rect 15565 15555 15623 15561
rect 15565 15521 15577 15555
rect 15611 15521 15623 15555
rect 15565 15515 15623 15521
rect 14918 15444 14924 15496
rect 14976 15484 14982 15496
rect 15105 15487 15163 15493
rect 15105 15484 15117 15487
rect 14976 15456 15117 15484
rect 14976 15444 14982 15456
rect 15105 15453 15117 15456
rect 15151 15453 15163 15487
rect 15212 15484 15240 15512
rect 15580 15484 15608 15515
rect 15856 15493 15884 15592
rect 21542 15580 21548 15632
rect 21600 15620 21606 15632
rect 21600 15592 22232 15620
rect 21600 15580 21606 15592
rect 18506 15561 18512 15564
rect 18500 15552 18512 15561
rect 18467 15524 18512 15552
rect 18500 15515 18512 15524
rect 18506 15512 18512 15515
rect 18564 15512 18570 15564
rect 21082 15512 21088 15564
rect 21140 15552 21146 15564
rect 21729 15555 21787 15561
rect 21729 15552 21741 15555
rect 21140 15524 21741 15552
rect 21140 15512 21146 15524
rect 21729 15521 21741 15524
rect 21775 15552 21787 15555
rect 22002 15552 22008 15564
rect 21775 15524 22008 15552
rect 21775 15521 21787 15524
rect 21729 15515 21787 15521
rect 22002 15512 22008 15524
rect 22060 15512 22066 15564
rect 22204 15561 22232 15592
rect 22189 15555 22247 15561
rect 22189 15521 22201 15555
rect 22235 15521 22247 15555
rect 22189 15515 22247 15521
rect 15212 15456 15608 15484
rect 15841 15487 15899 15493
rect 15105 15447 15163 15453
rect 15841 15453 15853 15487
rect 15887 15453 15899 15487
rect 15841 15447 15899 15453
rect 13372 15388 14320 15416
rect 4157 15351 4215 15357
rect 4157 15317 4169 15351
rect 4203 15348 4215 15351
rect 4246 15348 4252 15360
rect 4203 15320 4252 15348
rect 4203 15317 4215 15320
rect 4157 15311 4215 15317
rect 4246 15308 4252 15320
rect 4304 15308 4310 15360
rect 8573 15351 8631 15357
rect 8573 15317 8585 15351
rect 8619 15348 8631 15351
rect 8754 15348 8760 15360
rect 8619 15320 8760 15348
rect 8619 15317 8631 15320
rect 8573 15311 8631 15317
rect 8754 15308 8760 15320
rect 8812 15308 8818 15360
rect 15120 15348 15148 15447
rect 18230 15444 18236 15496
rect 18288 15444 18294 15496
rect 21818 15444 21824 15496
rect 21876 15444 21882 15496
rect 22281 15487 22339 15493
rect 22281 15484 22293 15487
rect 21928 15456 22293 15484
rect 15473 15419 15531 15425
rect 15473 15385 15485 15419
rect 15519 15416 15531 15419
rect 15930 15416 15936 15428
rect 15519 15388 15936 15416
rect 15519 15385 15531 15388
rect 15473 15379 15531 15385
rect 15930 15376 15936 15388
rect 15988 15376 15994 15428
rect 21450 15376 21456 15428
rect 21508 15416 21514 15428
rect 21928 15416 21956 15456
rect 22281 15453 22293 15456
rect 22327 15453 22339 15487
rect 22281 15447 22339 15453
rect 21508 15388 21956 15416
rect 22097 15419 22155 15425
rect 21508 15376 21514 15388
rect 22097 15385 22109 15419
rect 22143 15416 22155 15419
rect 22462 15416 22468 15428
rect 22143 15388 22468 15416
rect 22143 15385 22155 15388
rect 22097 15379 22155 15385
rect 22462 15376 22468 15388
rect 22520 15376 22526 15428
rect 15654 15348 15660 15360
rect 15120 15320 15660 15348
rect 15654 15308 15660 15320
rect 15712 15308 15718 15360
rect 15746 15308 15752 15360
rect 15804 15308 15810 15360
rect 19426 15308 19432 15360
rect 19484 15348 19490 15360
rect 19613 15351 19671 15357
rect 19613 15348 19625 15351
rect 19484 15320 19625 15348
rect 19484 15308 19490 15320
rect 19613 15317 19625 15320
rect 19659 15317 19671 15351
rect 19613 15311 19671 15317
rect 22278 15308 22284 15360
rect 22336 15308 22342 15360
rect 552 15258 23368 15280
rect 552 15206 3662 15258
rect 3714 15206 3726 15258
rect 3778 15206 3790 15258
rect 3842 15206 3854 15258
rect 3906 15206 3918 15258
rect 3970 15206 23368 15258
rect 552 15184 23368 15206
rect 5997 15147 6055 15153
rect 5997 15113 6009 15147
rect 6043 15144 6055 15147
rect 11238 15144 11244 15156
rect 6043 15116 11244 15144
rect 6043 15113 6055 15116
rect 5997 15107 6055 15113
rect 11238 15104 11244 15116
rect 11296 15104 11302 15156
rect 13814 15104 13820 15156
rect 13872 15144 13878 15156
rect 13909 15147 13967 15153
rect 13909 15144 13921 15147
rect 13872 15116 13921 15144
rect 13872 15104 13878 15116
rect 13909 15113 13921 15116
rect 13955 15113 13967 15147
rect 13909 15107 13967 15113
rect 16022 15104 16028 15156
rect 16080 15144 16086 15156
rect 17954 15144 17960 15156
rect 16080 15116 17960 15144
rect 16080 15104 16086 15116
rect 17954 15104 17960 15116
rect 18012 15144 18018 15156
rect 18012 15116 18368 15144
rect 18012 15104 18018 15116
rect 4525 15079 4583 15085
rect 4525 15045 4537 15079
rect 4571 15076 4583 15079
rect 4571 15048 5856 15076
rect 4571 15045 4583 15048
rect 4525 15039 4583 15045
rect 4246 14968 4252 15020
rect 4304 14968 4310 15020
rect 4706 14968 4712 15020
rect 4764 14968 4770 15020
rect 5828 15017 5856 15048
rect 10962 15036 10968 15088
rect 11020 15036 11026 15088
rect 16482 15036 16488 15088
rect 16540 15076 16546 15088
rect 16577 15079 16635 15085
rect 16577 15076 16589 15079
rect 16540 15048 16589 15076
rect 16540 15036 16546 15048
rect 16577 15045 16589 15048
rect 16623 15045 16635 15079
rect 16577 15039 16635 15045
rect 5813 15011 5871 15017
rect 5813 14977 5825 15011
rect 5859 15008 5871 15011
rect 5902 15008 5908 15020
rect 5859 14980 5908 15008
rect 5859 14977 5871 14980
rect 5813 14971 5871 14977
rect 5902 14968 5908 14980
rect 5960 14968 5966 15020
rect 10873 15011 10931 15017
rect 10873 14977 10885 15011
rect 10919 15008 10931 15011
rect 10980 15008 11008 15036
rect 10919 14980 11008 15008
rect 10919 14977 10931 14980
rect 10873 14971 10931 14977
rect 15746 14968 15752 15020
rect 15804 15008 15810 15020
rect 16209 15011 16267 15017
rect 16209 15008 16221 15011
rect 15804 14980 16221 15008
rect 15804 14968 15810 14980
rect 16209 14977 16221 14980
rect 16255 15008 16267 15011
rect 16255 14980 16896 15008
rect 16255 14977 16267 14980
rect 16209 14971 16267 14977
rect 4154 14900 4160 14952
rect 4212 14900 4218 14952
rect 4801 14943 4859 14949
rect 4801 14909 4813 14943
rect 4847 14940 4859 14943
rect 4982 14940 4988 14952
rect 4847 14912 4988 14940
rect 4847 14909 4859 14912
rect 4801 14903 4859 14909
rect 4982 14900 4988 14912
rect 5040 14900 5046 14952
rect 5721 14943 5779 14949
rect 5721 14909 5733 14943
rect 5767 14940 5779 14943
rect 7006 14940 7012 14952
rect 5767 14912 7012 14940
rect 5767 14909 5779 14912
rect 5721 14903 5779 14909
rect 7006 14900 7012 14912
rect 7064 14900 7070 14952
rect 10965 14943 11023 14949
rect 10965 14909 10977 14943
rect 11011 14940 11023 14943
rect 11054 14940 11060 14952
rect 11011 14912 11060 14940
rect 11011 14909 11023 14912
rect 10965 14903 11023 14909
rect 11054 14900 11060 14912
rect 11112 14900 11118 14952
rect 12618 14900 12624 14952
rect 12676 14900 12682 14952
rect 13081 14943 13139 14949
rect 13081 14909 13093 14943
rect 13127 14940 13139 14943
rect 13725 14943 13783 14949
rect 13725 14940 13737 14943
rect 13127 14912 13737 14940
rect 13127 14909 13139 14912
rect 13081 14903 13139 14909
rect 13725 14909 13737 14912
rect 13771 14940 13783 14943
rect 14182 14940 14188 14952
rect 13771 14912 14188 14940
rect 13771 14909 13783 14912
rect 13725 14903 13783 14909
rect 14182 14900 14188 14912
rect 14240 14900 14246 14952
rect 15470 14900 15476 14952
rect 15528 14940 15534 14952
rect 16022 14940 16028 14952
rect 15528 14912 16028 14940
rect 15528 14900 15534 14912
rect 16022 14900 16028 14912
rect 16080 14900 16086 14952
rect 16117 14943 16175 14949
rect 16117 14909 16129 14943
rect 16163 14909 16175 14943
rect 16117 14903 16175 14909
rect 16301 14943 16359 14949
rect 16301 14909 16313 14943
rect 16347 14940 16359 14943
rect 16574 14940 16580 14952
rect 16347 14912 16580 14940
rect 16347 14909 16359 14912
rect 16301 14903 16359 14909
rect 12636 14872 12664 14900
rect 13541 14875 13599 14881
rect 13541 14872 13553 14875
rect 12636 14844 13553 14872
rect 13541 14841 13553 14844
rect 13587 14841 13599 14875
rect 16132 14872 16160 14903
rect 16574 14900 16580 14912
rect 16632 14900 16638 14952
rect 16758 14900 16764 14952
rect 16816 14900 16822 14952
rect 16868 14949 16896 14980
rect 16853 14943 16911 14949
rect 16853 14909 16865 14943
rect 16899 14909 16911 14943
rect 18340 14940 18368 15116
rect 18414 15104 18420 15156
rect 18472 15144 18478 15156
rect 18785 15147 18843 15153
rect 18785 15144 18797 15147
rect 18472 15116 18797 15144
rect 18472 15104 18478 15116
rect 18785 15113 18797 15116
rect 18831 15113 18843 15147
rect 18785 15107 18843 15113
rect 21542 15104 21548 15156
rect 21600 15104 21606 15156
rect 21560 15076 21588 15104
rect 21284 15048 21588 15076
rect 20257 15011 20315 15017
rect 20257 14977 20269 15011
rect 20303 15008 20315 15011
rect 20346 15008 20352 15020
rect 20303 14980 20352 15008
rect 20303 14977 20315 14980
rect 20257 14971 20315 14977
rect 20346 14968 20352 14980
rect 20404 15008 20410 15020
rect 20898 15008 20904 15020
rect 20404 14980 20904 15008
rect 20404 14968 20410 14980
rect 20898 14968 20904 14980
rect 20956 15008 20962 15020
rect 21284 15017 21312 15048
rect 21269 15011 21327 15017
rect 21269 15008 21281 15011
rect 20956 14980 21281 15008
rect 20956 14968 20962 14980
rect 21269 14977 21281 14980
rect 21315 14977 21327 15011
rect 21269 14971 21327 14977
rect 21450 14968 21456 15020
rect 21508 15008 21514 15020
rect 21545 15011 21603 15017
rect 21545 15008 21557 15011
rect 21508 14980 21557 15008
rect 21508 14968 21514 14980
rect 21545 14977 21557 14980
rect 21591 14977 21603 15011
rect 21545 14971 21603 14977
rect 18693 14943 18751 14949
rect 18693 14940 18705 14943
rect 18340 14912 18705 14940
rect 16853 14903 16911 14909
rect 18693 14909 18705 14912
rect 18739 14909 18751 14943
rect 18693 14903 18751 14909
rect 18877 14943 18935 14949
rect 18877 14909 18889 14943
rect 18923 14940 18935 14943
rect 19426 14940 19432 14952
rect 18923 14912 19432 14940
rect 18923 14909 18935 14912
rect 18877 14903 18935 14909
rect 19426 14900 19432 14912
rect 19484 14900 19490 14952
rect 21177 14943 21235 14949
rect 21177 14909 21189 14943
rect 21223 14940 21235 14943
rect 21358 14940 21364 14952
rect 21223 14912 21364 14940
rect 21223 14909 21235 14912
rect 21177 14903 21235 14909
rect 21358 14900 21364 14912
rect 21416 14900 21422 14952
rect 22002 14900 22008 14952
rect 22060 14900 22066 14952
rect 16776 14872 16804 14900
rect 16132 14844 16804 14872
rect 13541 14835 13599 14841
rect 19886 14832 19892 14884
rect 19944 14832 19950 14884
rect 20070 14832 20076 14884
rect 20128 14872 20134 14884
rect 20622 14872 20628 14884
rect 20128 14844 20628 14872
rect 20128 14832 20134 14844
rect 20622 14832 20628 14844
rect 20680 14832 20686 14884
rect 21818 14832 21824 14884
rect 21876 14832 21882 14884
rect 22189 14875 22247 14881
rect 22189 14841 22201 14875
rect 22235 14872 22247 14875
rect 22554 14872 22560 14884
rect 22235 14844 22560 14872
rect 22235 14841 22247 14844
rect 22189 14835 22247 14841
rect 22554 14832 22560 14844
rect 22612 14872 22618 14884
rect 22830 14872 22836 14884
rect 22612 14844 22836 14872
rect 22612 14832 22618 14844
rect 22830 14832 22836 14844
rect 22888 14832 22894 14884
rect 5166 14764 5172 14816
rect 5224 14764 5230 14816
rect 5350 14764 5356 14816
rect 5408 14764 5414 14816
rect 11333 14807 11391 14813
rect 11333 14773 11345 14807
rect 11379 14804 11391 14807
rect 11514 14804 11520 14816
rect 11379 14776 11520 14804
rect 11379 14773 11391 14776
rect 11333 14767 11391 14773
rect 11514 14764 11520 14776
rect 11572 14764 11578 14816
rect 12253 14807 12311 14813
rect 12253 14773 12265 14807
rect 12299 14804 12311 14807
rect 12802 14804 12808 14816
rect 12299 14776 12808 14804
rect 12299 14773 12311 14776
rect 12253 14767 12311 14773
rect 12802 14764 12808 14776
rect 12860 14764 12866 14816
rect 16390 14764 16396 14816
rect 16448 14804 16454 14816
rect 16485 14807 16543 14813
rect 16485 14804 16497 14807
rect 16448 14776 16497 14804
rect 16448 14764 16454 14776
rect 16485 14773 16497 14776
rect 16531 14773 16543 14807
rect 16485 14767 16543 14773
rect 552 14714 23368 14736
rect 552 14662 4322 14714
rect 4374 14662 4386 14714
rect 4438 14662 4450 14714
rect 4502 14662 4514 14714
rect 4566 14662 4578 14714
rect 4630 14662 23368 14714
rect 552 14640 23368 14662
rect 2958 14560 2964 14612
rect 3016 14600 3022 14612
rect 3053 14603 3111 14609
rect 3053 14600 3065 14603
rect 3016 14572 3065 14600
rect 3016 14560 3022 14572
rect 3053 14569 3065 14572
rect 3099 14600 3111 14603
rect 3418 14600 3424 14612
rect 3099 14572 3424 14600
rect 3099 14569 3111 14572
rect 3053 14563 3111 14569
rect 3418 14560 3424 14572
rect 3476 14560 3482 14612
rect 4525 14603 4583 14609
rect 4525 14569 4537 14603
rect 4571 14600 4583 14603
rect 5350 14600 5356 14612
rect 4571 14572 5356 14600
rect 4571 14569 4583 14572
rect 4525 14563 4583 14569
rect 5350 14560 5356 14572
rect 5408 14560 5414 14612
rect 19334 14600 19340 14612
rect 17604 14572 19340 14600
rect 4154 14492 4160 14544
rect 4212 14532 4218 14544
rect 10042 14532 10048 14544
rect 4212 14504 4568 14532
rect 4212 14492 4218 14504
rect 2685 14467 2743 14473
rect 2685 14433 2697 14467
rect 2731 14464 2743 14467
rect 2774 14464 2780 14476
rect 2731 14436 2780 14464
rect 2731 14433 2743 14436
rect 2685 14427 2743 14433
rect 2774 14424 2780 14436
rect 2832 14424 2838 14476
rect 2866 14424 2872 14476
rect 2924 14424 2930 14476
rect 4246 14424 4252 14476
rect 4304 14464 4310 14476
rect 4540 14473 4568 14504
rect 9232 14504 10048 14532
rect 4341 14467 4399 14473
rect 4341 14464 4353 14467
rect 4304 14436 4353 14464
rect 4304 14424 4310 14436
rect 4341 14433 4353 14436
rect 4387 14433 4399 14467
rect 4341 14427 4399 14433
rect 4525 14467 4583 14473
rect 4525 14433 4537 14467
rect 4571 14433 4583 14467
rect 4525 14427 4583 14433
rect 5166 14424 5172 14476
rect 5224 14424 5230 14476
rect 5997 14467 6055 14473
rect 5997 14433 6009 14467
rect 6043 14464 6055 14467
rect 6086 14464 6092 14476
rect 6043 14436 6092 14464
rect 6043 14433 6055 14436
rect 5997 14427 6055 14433
rect 6086 14424 6092 14436
rect 6144 14464 6150 14476
rect 7190 14464 7196 14476
rect 6144 14436 7196 14464
rect 6144 14424 6150 14436
rect 7190 14424 7196 14436
rect 7248 14424 7254 14476
rect 8018 14424 8024 14476
rect 8076 14424 8082 14476
rect 9030 14424 9036 14476
rect 9088 14464 9094 14476
rect 9232 14473 9260 14504
rect 10042 14492 10048 14504
rect 10100 14492 10106 14544
rect 15746 14492 15752 14544
rect 15804 14492 15810 14544
rect 9217 14467 9275 14473
rect 9217 14464 9229 14467
rect 9088 14436 9229 14464
rect 9088 14424 9094 14436
rect 9217 14433 9229 14436
rect 9263 14433 9275 14467
rect 9217 14427 9275 14433
rect 9310 14467 9368 14473
rect 9310 14433 9322 14467
rect 9356 14433 9368 14467
rect 9310 14427 9368 14433
rect 5261 14399 5319 14405
rect 5261 14365 5273 14399
rect 5307 14396 5319 14399
rect 5442 14396 5448 14408
rect 5307 14368 5448 14396
rect 5307 14365 5319 14368
rect 5261 14359 5319 14365
rect 5442 14356 5448 14368
rect 5500 14356 5506 14408
rect 5902 14356 5908 14408
rect 5960 14356 5966 14408
rect 8113 14399 8171 14405
rect 8113 14365 8125 14399
rect 8159 14396 8171 14399
rect 8386 14396 8392 14408
rect 8159 14368 8392 14396
rect 8159 14365 8171 14368
rect 8113 14359 8171 14365
rect 8386 14356 8392 14368
rect 8444 14356 8450 14408
rect 9324 14396 9352 14427
rect 15470 14424 15476 14476
rect 15528 14464 15534 14476
rect 15565 14467 15623 14473
rect 15565 14464 15577 14467
rect 15528 14436 15577 14464
rect 15528 14424 15534 14436
rect 15565 14433 15577 14436
rect 15611 14433 15623 14467
rect 15565 14427 15623 14433
rect 15654 14424 15660 14476
rect 15712 14424 15718 14476
rect 15930 14424 15936 14476
rect 15988 14424 15994 14476
rect 16117 14467 16175 14473
rect 16117 14433 16129 14467
rect 16163 14433 16175 14467
rect 16117 14427 16175 14433
rect 8956 14368 9352 14396
rect 16132 14396 16160 14427
rect 16390 14424 16396 14476
rect 16448 14424 16454 14476
rect 16482 14424 16488 14476
rect 16540 14424 16546 14476
rect 17494 14396 17500 14408
rect 16132 14368 17500 14396
rect 5537 14331 5595 14337
rect 5537 14297 5549 14331
rect 5583 14328 5595 14331
rect 5994 14328 6000 14340
rect 5583 14300 6000 14328
rect 5583 14297 5595 14300
rect 5537 14291 5595 14297
rect 5994 14288 6000 14300
rect 6052 14288 6058 14340
rect 8956 14272 8984 14368
rect 17494 14356 17500 14368
rect 17552 14356 17558 14408
rect 9585 14331 9643 14337
rect 9585 14297 9597 14331
rect 9631 14328 9643 14331
rect 9674 14328 9680 14340
rect 9631 14300 9680 14328
rect 9631 14297 9643 14300
rect 9585 14291 9643 14297
rect 9674 14288 9680 14300
rect 9732 14288 9738 14340
rect 15010 14288 15016 14340
rect 15068 14328 15074 14340
rect 16209 14331 16267 14337
rect 16209 14328 16221 14331
rect 15068 14300 16221 14328
rect 15068 14288 15074 14300
rect 16209 14297 16221 14300
rect 16255 14328 16267 14331
rect 17604 14328 17632 14572
rect 19334 14560 19340 14572
rect 19392 14560 19398 14612
rect 21082 14600 21088 14612
rect 20180 14572 21088 14600
rect 19705 14535 19763 14541
rect 18984 14504 19564 14532
rect 17770 14424 17776 14476
rect 17828 14464 17834 14476
rect 18984 14473 19012 14504
rect 18969 14467 19027 14473
rect 18969 14464 18981 14467
rect 17828 14436 18981 14464
rect 17828 14424 17834 14436
rect 18969 14433 18981 14436
rect 19015 14433 19027 14467
rect 18969 14427 19027 14433
rect 19153 14467 19211 14473
rect 19153 14433 19165 14467
rect 19199 14464 19211 14467
rect 19426 14464 19432 14476
rect 19199 14436 19432 14464
rect 19199 14433 19211 14436
rect 19153 14427 19211 14433
rect 19426 14424 19432 14436
rect 19484 14424 19490 14476
rect 19536 14473 19564 14504
rect 19705 14501 19717 14535
rect 19751 14501 19763 14535
rect 19705 14495 19763 14501
rect 19521 14467 19579 14473
rect 19521 14433 19533 14467
rect 19567 14433 19579 14467
rect 19720 14464 19748 14495
rect 19797 14467 19855 14473
rect 19797 14464 19809 14467
rect 19720 14436 19809 14464
rect 19521 14427 19579 14433
rect 19797 14433 19809 14436
rect 19843 14433 19855 14467
rect 19797 14427 19855 14433
rect 19886 14424 19892 14476
rect 19944 14464 19950 14476
rect 20180 14473 20208 14572
rect 21082 14560 21088 14572
rect 21140 14560 21146 14612
rect 20272 14504 20576 14532
rect 19981 14467 20039 14473
rect 19981 14464 19993 14467
rect 19944 14436 19993 14464
rect 19944 14424 19950 14436
rect 19981 14433 19993 14436
rect 20027 14433 20039 14467
rect 19981 14427 20039 14433
rect 20165 14467 20223 14473
rect 20165 14433 20177 14467
rect 20211 14433 20223 14467
rect 20165 14427 20223 14433
rect 19242 14356 19248 14408
rect 19300 14396 19306 14408
rect 19705 14399 19763 14405
rect 19705 14396 19717 14399
rect 19300 14368 19717 14396
rect 19300 14356 19306 14368
rect 19705 14365 19717 14368
rect 19751 14365 19763 14399
rect 19705 14359 19763 14365
rect 19996 14396 20024 14427
rect 20272 14396 20300 14504
rect 20346 14424 20352 14476
rect 20404 14424 20410 14476
rect 20548 14473 20576 14504
rect 20441 14467 20499 14473
rect 20441 14433 20453 14467
rect 20487 14433 20499 14467
rect 20441 14427 20499 14433
rect 20533 14467 20591 14473
rect 20533 14433 20545 14467
rect 20579 14433 20591 14467
rect 20533 14427 20591 14433
rect 19996 14368 20300 14396
rect 20456 14396 20484 14427
rect 20622 14424 20628 14476
rect 20680 14464 20686 14476
rect 20717 14467 20775 14473
rect 20717 14464 20729 14467
rect 20680 14436 20729 14464
rect 20680 14424 20686 14436
rect 20717 14433 20729 14436
rect 20763 14433 20775 14467
rect 20717 14427 20775 14433
rect 20456 14368 20668 14396
rect 16255 14300 17632 14328
rect 16255 14297 16267 14300
rect 16209 14291 16267 14297
rect 6273 14263 6331 14269
rect 6273 14229 6285 14263
rect 6319 14260 6331 14263
rect 6730 14260 6736 14272
rect 6319 14232 6736 14260
rect 6319 14229 6331 14232
rect 6273 14223 6331 14229
rect 6730 14220 6736 14232
rect 6788 14220 6794 14272
rect 8297 14263 8355 14269
rect 8297 14229 8309 14263
rect 8343 14260 8355 14263
rect 8938 14260 8944 14272
rect 8343 14232 8944 14260
rect 8343 14229 8355 14232
rect 8297 14223 8355 14229
rect 8938 14220 8944 14232
rect 8996 14220 9002 14272
rect 15378 14220 15384 14272
rect 15436 14220 15442 14272
rect 16669 14263 16727 14269
rect 16669 14229 16681 14263
rect 16715 14260 16727 14263
rect 16850 14260 16856 14272
rect 16715 14232 16856 14260
rect 16715 14229 16727 14232
rect 16669 14223 16727 14229
rect 16850 14220 16856 14232
rect 16908 14220 16914 14272
rect 19153 14263 19211 14269
rect 19153 14229 19165 14263
rect 19199 14260 19211 14263
rect 19260 14260 19288 14356
rect 19337 14331 19395 14337
rect 19337 14297 19349 14331
rect 19383 14328 19395 14331
rect 19996 14328 20024 14368
rect 19383 14300 20024 14328
rect 19383 14297 19395 14300
rect 19337 14291 19395 14297
rect 19199 14232 19288 14260
rect 19199 14229 19211 14232
rect 19153 14223 19211 14229
rect 19610 14220 19616 14272
rect 19668 14260 19674 14272
rect 19889 14263 19947 14269
rect 19889 14260 19901 14263
rect 19668 14232 19901 14260
rect 19668 14220 19674 14232
rect 19889 14229 19901 14232
rect 19935 14229 19947 14263
rect 19889 14223 19947 14229
rect 20162 14220 20168 14272
rect 20220 14220 20226 14272
rect 20640 14269 20668 14368
rect 20625 14263 20683 14269
rect 20625 14229 20637 14263
rect 20671 14260 20683 14263
rect 20806 14260 20812 14272
rect 20671 14232 20812 14260
rect 20671 14229 20683 14232
rect 20625 14223 20683 14229
rect 20806 14220 20812 14232
rect 20864 14220 20870 14272
rect 552 14170 23368 14192
rect 552 14118 3662 14170
rect 3714 14118 3726 14170
rect 3778 14118 3790 14170
rect 3842 14118 3854 14170
rect 3906 14118 3918 14170
rect 3970 14118 23368 14170
rect 552 14096 23368 14118
rect 7009 14059 7067 14065
rect 7009 14025 7021 14059
rect 7055 14056 7067 14059
rect 8021 14059 8079 14065
rect 7055 14028 7880 14056
rect 7055 14025 7067 14028
rect 7009 14019 7067 14025
rect 3053 13991 3111 13997
rect 3053 13957 3065 13991
rect 3099 13957 3111 13991
rect 3053 13951 3111 13957
rect 2774 13812 2780 13864
rect 2832 13812 2838 13864
rect 2866 13812 2872 13864
rect 2924 13812 2930 13864
rect 3068 13852 3096 13951
rect 5166 13948 5172 14000
rect 5224 13988 5230 14000
rect 5537 13991 5595 13997
rect 5537 13988 5549 13991
rect 5224 13960 5549 13988
rect 5224 13948 5230 13960
rect 5537 13957 5549 13960
rect 5583 13957 5595 13991
rect 5537 13951 5595 13957
rect 6457 13991 6515 13997
rect 6457 13957 6469 13991
rect 6503 13988 6515 13991
rect 6503 13960 7512 13988
rect 6503 13957 6515 13960
rect 6457 13951 6515 13957
rect 3142 13880 3148 13932
rect 3200 13920 3206 13932
rect 5261 13923 5319 13929
rect 3200 13892 3648 13920
rect 3200 13880 3206 13892
rect 3237 13855 3295 13861
rect 3237 13852 3249 13855
rect 3068 13824 3249 13852
rect 3237 13821 3249 13824
rect 3283 13821 3295 13855
rect 3237 13815 3295 13821
rect 3418 13812 3424 13864
rect 3476 13812 3482 13864
rect 3620 13861 3648 13892
rect 5261 13889 5273 13923
rect 5307 13920 5319 13923
rect 5442 13920 5448 13932
rect 5307 13892 5448 13920
rect 5307 13889 5319 13892
rect 5261 13883 5319 13889
rect 5442 13880 5448 13892
rect 5500 13880 5506 13932
rect 5994 13880 6000 13932
rect 6052 13880 6058 13932
rect 6638 13880 6644 13932
rect 6696 13880 6702 13932
rect 6748 13892 7328 13920
rect 6748 13864 6776 13892
rect 3605 13855 3663 13861
rect 3605 13821 3617 13855
rect 3651 13821 3663 13855
rect 3605 13815 3663 13821
rect 6086 13812 6092 13864
rect 6144 13812 6150 13864
rect 6730 13812 6736 13864
rect 6788 13812 6794 13864
rect 7300 13861 7328 13892
rect 7193 13855 7251 13861
rect 7193 13852 7205 13855
rect 6840 13824 7205 13852
rect 3053 13787 3111 13793
rect 3053 13753 3065 13787
rect 3099 13784 3111 13787
rect 3142 13784 3148 13796
rect 3099 13756 3148 13784
rect 3099 13753 3111 13756
rect 3053 13747 3111 13753
rect 3142 13744 3148 13756
rect 3200 13744 3206 13796
rect 3510 13744 3516 13796
rect 3568 13744 3574 13796
rect 6638 13744 6644 13796
rect 6696 13784 6702 13796
rect 6840 13784 6868 13824
rect 7193 13821 7205 13824
rect 7239 13821 7251 13855
rect 7193 13815 7251 13821
rect 7286 13855 7344 13861
rect 7286 13821 7298 13855
rect 7332 13821 7344 13855
rect 7484 13852 7512 13960
rect 7852 13920 7880 14028
rect 8021 14025 8033 14059
rect 8067 14056 8079 14059
rect 9490 14056 9496 14068
rect 8067 14028 9496 14056
rect 8067 14025 8079 14028
rect 8021 14019 8079 14025
rect 9490 14016 9496 14028
rect 9548 14016 9554 14068
rect 10689 14059 10747 14065
rect 10689 14025 10701 14059
rect 10735 14056 10747 14059
rect 11238 14056 11244 14068
rect 10735 14028 11244 14056
rect 10735 14025 10747 14028
rect 10689 14019 10747 14025
rect 11238 14016 11244 14028
rect 11296 14056 11302 14068
rect 11977 14059 12035 14065
rect 11977 14056 11989 14059
rect 11296 14028 11989 14056
rect 11296 14016 11302 14028
rect 11977 14025 11989 14028
rect 12023 14025 12035 14059
rect 11977 14019 12035 14025
rect 13906 14016 13912 14068
rect 13964 14056 13970 14068
rect 14093 14059 14151 14065
rect 14093 14056 14105 14059
rect 13964 14028 14105 14056
rect 13964 14016 13970 14028
rect 14093 14025 14105 14028
rect 14139 14025 14151 14059
rect 14093 14019 14151 14025
rect 15654 14016 15660 14068
rect 15712 14056 15718 14068
rect 16206 14056 16212 14068
rect 15712 14028 16212 14056
rect 15712 14016 15718 14028
rect 16206 14016 16212 14028
rect 16264 14056 16270 14068
rect 16669 14059 16727 14065
rect 16669 14056 16681 14059
rect 16264 14028 16681 14056
rect 16264 14016 16270 14028
rect 16669 14025 16681 14028
rect 16715 14025 16727 14059
rect 16669 14019 16727 14025
rect 17494 14016 17500 14068
rect 17552 14056 17558 14068
rect 18141 14059 18199 14065
rect 18141 14056 18153 14059
rect 17552 14028 18153 14056
rect 17552 14016 17558 14028
rect 18141 14025 18153 14028
rect 18187 14025 18199 14059
rect 18141 14019 18199 14025
rect 20162 14016 20168 14068
rect 20220 14016 20226 14068
rect 20625 14059 20683 14065
rect 20625 14025 20637 14059
rect 20671 14056 20683 14059
rect 20671 14028 20852 14056
rect 20671 14025 20683 14028
rect 20625 14019 20683 14025
rect 8846 13948 8852 14000
rect 8904 13988 8910 14000
rect 8904 13960 11376 13988
rect 8904 13948 8910 13960
rect 7852 13892 8892 13920
rect 8018 13852 8024 13864
rect 8076 13861 8082 13864
rect 8076 13855 8109 13861
rect 7484 13824 8024 13852
rect 7286 13815 7344 13821
rect 8018 13812 8024 13824
rect 8097 13821 8109 13855
rect 8076 13815 8109 13821
rect 8205 13855 8263 13861
rect 8205 13821 8217 13855
rect 8251 13852 8263 13855
rect 8386 13852 8392 13864
rect 8251 13824 8392 13852
rect 8251 13821 8263 13824
rect 8205 13815 8263 13821
rect 8076 13812 8082 13815
rect 8386 13812 8392 13824
rect 8444 13812 8450 13864
rect 8864 13852 8892 13892
rect 8938 13880 8944 13932
rect 8996 13880 9002 13932
rect 9769 13923 9827 13929
rect 9769 13920 9781 13923
rect 9140 13892 9781 13920
rect 8864 13824 8984 13852
rect 6696 13756 6868 13784
rect 7561 13787 7619 13793
rect 6696 13744 6702 13756
rect 7561 13753 7573 13787
rect 7607 13784 7619 13787
rect 8846 13784 8852 13796
rect 7607 13756 8852 13784
rect 7607 13753 7619 13756
rect 7561 13747 7619 13753
rect 8846 13744 8852 13756
rect 8904 13744 8910 13796
rect 8956 13784 8984 13824
rect 9030 13812 9036 13864
rect 9088 13812 9094 13864
rect 9140 13784 9168 13892
rect 9769 13889 9781 13892
rect 9815 13889 9827 13923
rect 9769 13883 9827 13889
rect 9677 13855 9735 13861
rect 9677 13821 9689 13855
rect 9723 13821 9735 13855
rect 9784 13852 9812 13883
rect 10597 13855 10655 13861
rect 10597 13852 10609 13855
rect 9784 13824 10609 13852
rect 9677 13815 9735 13821
rect 10597 13821 10609 13824
rect 10643 13821 10655 13855
rect 10781 13855 10839 13861
rect 10781 13852 10793 13855
rect 10597 13815 10655 13821
rect 10704 13824 10793 13852
rect 8956 13756 9168 13784
rect 9692 13784 9720 13815
rect 10704 13784 10732 13824
rect 10781 13821 10793 13824
rect 10827 13852 10839 13855
rect 11054 13852 11060 13864
rect 10827 13824 11060 13852
rect 10827 13821 10839 13824
rect 10781 13815 10839 13821
rect 11054 13812 11060 13824
rect 11112 13812 11118 13864
rect 11238 13812 11244 13864
rect 11296 13812 11302 13864
rect 11348 13861 11376 13960
rect 17770 13948 17776 14000
rect 17828 13988 17834 14000
rect 20717 13991 20775 13997
rect 17828 13960 19012 13988
rect 17828 13948 17834 13960
rect 13262 13880 13268 13932
rect 13320 13920 13326 13932
rect 18230 13920 18236 13932
rect 13320 13892 13952 13920
rect 13320 13880 13326 13892
rect 11333 13855 11391 13861
rect 11333 13821 11345 13855
rect 11379 13821 11391 13855
rect 11333 13815 11391 13821
rect 9692 13756 10732 13784
rect 11348 13784 11376 13815
rect 11514 13812 11520 13864
rect 11572 13852 11578 13864
rect 11572 13824 12020 13852
rect 11572 13812 11578 13824
rect 11992 13793 12020 13824
rect 12894 13812 12900 13864
rect 12952 13852 12958 13864
rect 13541 13855 13599 13861
rect 13541 13852 13553 13855
rect 12952 13824 13553 13852
rect 12952 13812 12958 13824
rect 13541 13821 13553 13824
rect 13587 13821 13599 13855
rect 13541 13815 13599 13821
rect 13630 13812 13636 13864
rect 13688 13812 13694 13864
rect 13924 13861 13952 13892
rect 17788 13892 18236 13920
rect 13817 13855 13875 13861
rect 13817 13852 13829 13855
rect 13740 13824 13829 13852
rect 11793 13787 11851 13793
rect 11793 13784 11805 13787
rect 11348 13756 11805 13784
rect 11793 13753 11805 13756
rect 11839 13753 11851 13787
rect 11992 13787 12051 13793
rect 11992 13756 12005 13787
rect 11793 13747 11851 13753
rect 11993 13753 12005 13756
rect 12039 13753 12051 13787
rect 12342 13784 12348 13796
rect 11993 13747 12051 13753
rect 12084 13756 12348 13784
rect 3786 13676 3792 13728
rect 3844 13676 3850 13728
rect 5718 13676 5724 13728
rect 5776 13676 5782 13728
rect 8662 13676 8668 13728
rect 8720 13676 8726 13728
rect 10045 13719 10103 13725
rect 10045 13685 10057 13719
rect 10091 13716 10103 13719
rect 10226 13716 10232 13728
rect 10091 13688 10232 13716
rect 10091 13685 10103 13688
rect 10045 13679 10103 13685
rect 10226 13676 10232 13688
rect 10284 13676 10290 13728
rect 11701 13719 11759 13725
rect 11701 13685 11713 13719
rect 11747 13716 11759 13719
rect 12084 13716 12112 13756
rect 12342 13744 12348 13756
rect 12400 13784 12406 13796
rect 13740 13784 13768 13824
rect 13817 13821 13829 13824
rect 13863 13821 13875 13855
rect 13817 13815 13875 13821
rect 13909 13855 13967 13861
rect 13909 13821 13921 13855
rect 13955 13821 13967 13855
rect 13909 13815 13967 13821
rect 14550 13812 14556 13864
rect 14608 13852 14614 13864
rect 15289 13855 15347 13861
rect 15289 13852 15301 13855
rect 14608 13824 15301 13852
rect 14608 13812 14614 13824
rect 15289 13821 15301 13824
rect 15335 13821 15347 13855
rect 15289 13815 15347 13821
rect 12400 13756 13768 13784
rect 15304 13784 15332 13815
rect 15378 13812 15384 13864
rect 15436 13852 15442 13864
rect 15545 13855 15603 13861
rect 15545 13852 15557 13855
rect 15436 13824 15557 13852
rect 15436 13812 15442 13824
rect 15545 13821 15557 13824
rect 15591 13821 15603 13855
rect 16761 13855 16819 13861
rect 16761 13852 16773 13855
rect 15545 13815 15603 13821
rect 15672 13824 16773 13852
rect 15672 13784 15700 13824
rect 16761 13821 16773 13824
rect 16807 13821 16819 13855
rect 16761 13815 16819 13821
rect 15304 13756 15700 13784
rect 16776 13784 16804 13815
rect 16850 13812 16856 13864
rect 16908 13852 16914 13864
rect 17017 13855 17075 13861
rect 17017 13852 17029 13855
rect 16908 13824 17029 13852
rect 16908 13812 16914 13824
rect 17017 13821 17029 13824
rect 17063 13821 17075 13855
rect 17788 13852 17816 13892
rect 18230 13880 18236 13892
rect 18288 13880 18294 13932
rect 18506 13880 18512 13932
rect 18564 13920 18570 13932
rect 18984 13929 19012 13960
rect 20717 13957 20729 13991
rect 20763 13957 20775 13991
rect 20824 13988 20852 14028
rect 20898 14016 20904 14068
rect 20956 14016 20962 14068
rect 22002 14016 22008 14068
rect 22060 14056 22066 14068
rect 22649 14059 22707 14065
rect 22649 14056 22661 14059
rect 22060 14028 22661 14056
rect 22060 14016 22066 14028
rect 22649 14025 22661 14028
rect 22695 14025 22707 14059
rect 22649 14019 22707 14025
rect 21913 13991 21971 13997
rect 20824 13960 21680 13988
rect 20717 13951 20775 13957
rect 18693 13923 18751 13929
rect 18693 13920 18705 13923
rect 18564 13892 18705 13920
rect 18564 13880 18570 13892
rect 18693 13889 18705 13892
rect 18739 13889 18751 13923
rect 18693 13883 18751 13889
rect 18969 13923 19027 13929
rect 18969 13889 18981 13923
rect 19015 13889 19027 13923
rect 19426 13920 19432 13932
rect 18969 13883 19027 13889
rect 19076 13892 19432 13920
rect 19076 13861 19104 13892
rect 19426 13880 19432 13892
rect 19484 13880 19490 13932
rect 19610 13880 19616 13932
rect 19668 13880 19674 13932
rect 19889 13923 19947 13929
rect 19889 13889 19901 13923
rect 19935 13920 19947 13923
rect 20257 13923 20315 13929
rect 20257 13920 20269 13923
rect 19935 13892 20269 13920
rect 19935 13889 19947 13892
rect 19889 13883 19947 13889
rect 20257 13889 20269 13892
rect 20303 13889 20315 13923
rect 20257 13883 20315 13889
rect 17017 13815 17075 13821
rect 17144 13824 17816 13852
rect 19061 13855 19119 13861
rect 17144 13784 17172 13824
rect 19061 13821 19073 13855
rect 19107 13821 19119 13855
rect 19061 13815 19119 13821
rect 19334 13812 19340 13864
rect 19392 13852 19398 13864
rect 19521 13855 19579 13861
rect 19521 13852 19533 13855
rect 19392 13824 19533 13852
rect 19392 13812 19398 13824
rect 19521 13821 19533 13824
rect 19567 13821 19579 13855
rect 19521 13815 19579 13821
rect 20441 13855 20499 13861
rect 20441 13821 20453 13855
rect 20487 13852 20499 13855
rect 20732 13852 20760 13951
rect 21450 13880 21456 13932
rect 21508 13880 21514 13932
rect 20487 13824 20760 13852
rect 20487 13821 20499 13824
rect 20441 13815 20499 13821
rect 20806 13812 20812 13864
rect 20864 13827 20870 13864
rect 20864 13821 20913 13827
rect 20864 13812 20867 13821
rect 16776 13756 17172 13784
rect 12400 13744 12406 13756
rect 20162 13744 20168 13796
rect 20220 13744 20226 13796
rect 20824 13790 20867 13812
rect 20855 13787 20867 13790
rect 20901 13787 20913 13821
rect 21542 13812 21548 13864
rect 21600 13812 21606 13864
rect 21652 13852 21680 13960
rect 21913 13957 21925 13991
rect 21959 13988 21971 13991
rect 22189 13991 22247 13997
rect 22189 13988 22201 13991
rect 21959 13960 22201 13988
rect 21959 13957 21971 13960
rect 21913 13951 21971 13957
rect 22189 13957 22201 13960
rect 22235 13957 22247 13991
rect 22189 13951 22247 13957
rect 22005 13923 22063 13929
rect 22005 13889 22017 13923
rect 22051 13920 22063 13923
rect 22557 13923 22615 13929
rect 22557 13920 22569 13923
rect 22051 13892 22569 13920
rect 22051 13889 22063 13892
rect 22005 13883 22063 13889
rect 22557 13889 22569 13892
rect 22603 13889 22615 13923
rect 22557 13883 22615 13889
rect 22097 13855 22155 13861
rect 22097 13852 22109 13855
rect 21652 13824 22109 13852
rect 22097 13821 22109 13824
rect 22143 13821 22155 13855
rect 22097 13815 22155 13821
rect 22373 13855 22431 13861
rect 22373 13821 22385 13855
rect 22419 13821 22431 13855
rect 22373 13815 22431 13821
rect 20855 13781 20913 13787
rect 21082 13744 21088 13796
rect 21140 13744 21146 13796
rect 22388 13784 22416 13815
rect 22462 13812 22468 13864
rect 22520 13852 22526 13864
rect 22741 13855 22799 13861
rect 22741 13852 22753 13855
rect 22520 13824 22753 13852
rect 22520 13812 22526 13824
rect 22741 13821 22753 13824
rect 22787 13821 22799 13855
rect 22741 13815 22799 13821
rect 22833 13855 22891 13861
rect 22833 13821 22845 13855
rect 22879 13821 22891 13855
rect 22833 13815 22891 13821
rect 22554 13784 22560 13796
rect 22388 13756 22560 13784
rect 22554 13744 22560 13756
rect 22612 13784 22618 13796
rect 22848 13784 22876 13815
rect 22612 13756 22876 13784
rect 22612 13744 22618 13756
rect 11747 13688 12112 13716
rect 12161 13719 12219 13725
rect 11747 13685 11759 13688
rect 11701 13679 11759 13685
rect 12161 13685 12173 13719
rect 12207 13716 12219 13719
rect 12710 13716 12716 13728
rect 12207 13688 12716 13716
rect 12207 13685 12219 13688
rect 12161 13679 12219 13685
rect 12710 13676 12716 13688
rect 12768 13676 12774 13728
rect 20714 13676 20720 13728
rect 20772 13716 20778 13728
rect 21100 13716 21128 13744
rect 20772 13688 21128 13716
rect 20772 13676 20778 13688
rect 552 13626 23368 13648
rect 552 13574 4322 13626
rect 4374 13574 4386 13626
rect 4438 13574 4450 13626
rect 4502 13574 4514 13626
rect 4566 13574 4578 13626
rect 4630 13574 23368 13626
rect 552 13552 23368 13574
rect 10045 13515 10103 13521
rect 10045 13512 10057 13515
rect 9508 13484 10057 13512
rect 9508 13456 9536 13484
rect 10045 13481 10057 13484
rect 10091 13512 10103 13515
rect 10689 13515 10747 13521
rect 10689 13512 10701 13515
rect 10091 13484 10701 13512
rect 10091 13481 10103 13484
rect 10045 13475 10103 13481
rect 10689 13481 10701 13484
rect 10735 13481 10747 13515
rect 12529 13515 12587 13521
rect 12529 13512 12541 13515
rect 10689 13475 10747 13481
rect 12406 13484 12541 13512
rect 3786 13404 3792 13456
rect 3844 13444 3850 13456
rect 4074 13447 4132 13453
rect 4074 13444 4086 13447
rect 3844 13416 4086 13444
rect 3844 13404 3850 13416
rect 4074 13413 4086 13416
rect 4120 13413 4132 13447
rect 4074 13407 4132 13413
rect 5718 13404 5724 13456
rect 5776 13444 5782 13456
rect 6273 13447 6331 13453
rect 6273 13444 6285 13447
rect 5776 13416 6285 13444
rect 5776 13404 5782 13416
rect 6273 13413 6285 13416
rect 6319 13413 6331 13447
rect 6273 13407 6331 13413
rect 9490 13404 9496 13456
rect 9548 13404 9554 13456
rect 9709 13447 9767 13453
rect 9709 13413 9721 13447
rect 9755 13444 9767 13447
rect 12406 13444 12434 13484
rect 12529 13481 12541 13484
rect 12575 13481 12587 13515
rect 12529 13475 12587 13481
rect 12894 13472 12900 13524
rect 12952 13512 12958 13524
rect 12952 13484 13768 13512
rect 12952 13472 12958 13484
rect 13630 13444 13636 13456
rect 9755 13416 10272 13444
rect 9755 13413 9767 13416
rect 9709 13407 9767 13413
rect 10244 13388 10272 13416
rect 10888 13416 12434 13444
rect 12820 13416 13636 13444
rect 5994 13336 6000 13388
rect 6052 13336 6058 13388
rect 6089 13379 6147 13385
rect 6089 13345 6101 13379
rect 6135 13376 6147 13379
rect 7006 13376 7012 13388
rect 6135 13348 7012 13376
rect 6135 13345 6147 13348
rect 6089 13339 6147 13345
rect 7006 13336 7012 13348
rect 7064 13376 7070 13388
rect 8202 13376 8208 13388
rect 7064 13348 8208 13376
rect 7064 13336 7070 13348
rect 8202 13336 8208 13348
rect 8260 13336 8266 13388
rect 9953 13379 10011 13385
rect 9953 13376 9965 13379
rect 9692 13348 9965 13376
rect 9692 13320 9720 13348
rect 9953 13345 9965 13348
rect 9999 13345 10011 13379
rect 9953 13339 10011 13345
rect 4341 13311 4399 13317
rect 4341 13277 4353 13311
rect 4387 13308 4399 13311
rect 4706 13308 4712 13320
rect 4387 13280 4712 13308
rect 4387 13277 4399 13280
rect 4341 13271 4399 13277
rect 4706 13268 4712 13280
rect 4764 13268 4770 13320
rect 9674 13268 9680 13320
rect 9732 13268 9738 13320
rect 9968 13308 9996 13339
rect 10226 13336 10232 13388
rect 10284 13376 10290 13388
rect 10505 13379 10563 13385
rect 10505 13376 10517 13379
rect 10284 13348 10517 13376
rect 10284 13336 10290 13348
rect 10505 13345 10517 13348
rect 10551 13345 10563 13379
rect 10505 13339 10563 13345
rect 10781 13379 10839 13385
rect 10781 13345 10793 13379
rect 10827 13345 10839 13379
rect 10781 13339 10839 13345
rect 10796 13308 10824 13339
rect 9968 13280 10824 13308
rect 6273 13243 6331 13249
rect 6273 13209 6285 13243
rect 6319 13240 6331 13243
rect 6638 13240 6644 13252
rect 6319 13212 6644 13240
rect 6319 13209 6331 13212
rect 6273 13203 6331 13209
rect 6638 13200 6644 13212
rect 6696 13200 6702 13252
rect 9861 13243 9919 13249
rect 9861 13209 9873 13243
rect 9907 13240 9919 13243
rect 9950 13240 9956 13252
rect 9907 13212 9956 13240
rect 9907 13209 9919 13212
rect 9861 13203 9919 13209
rect 9950 13200 9956 13212
rect 10008 13240 10014 13252
rect 10888 13240 10916 13416
rect 12820 13388 12848 13416
rect 12342 13336 12348 13388
rect 12400 13376 12406 13388
rect 12437 13379 12495 13385
rect 12437 13376 12449 13379
rect 12400 13348 12449 13376
rect 12400 13336 12406 13348
rect 12437 13345 12449 13348
rect 12483 13345 12495 13379
rect 12437 13339 12495 13345
rect 12710 13336 12716 13388
rect 12768 13336 12774 13388
rect 12802 13336 12808 13388
rect 12860 13336 12866 13388
rect 12894 13336 12900 13388
rect 12952 13336 12958 13388
rect 13170 13336 13176 13388
rect 13228 13336 13234 13388
rect 13262 13336 13268 13388
rect 13320 13336 13326 13388
rect 13556 13385 13584 13416
rect 13630 13404 13636 13416
rect 13688 13404 13694 13456
rect 13740 13444 13768 13484
rect 13814 13472 13820 13524
rect 13872 13512 13878 13524
rect 14461 13515 14519 13521
rect 14461 13512 14473 13515
rect 13872 13484 14473 13512
rect 13872 13472 13878 13484
rect 14200 13453 14228 13484
rect 14461 13481 14473 13484
rect 14507 13481 14519 13515
rect 21910 13512 21916 13524
rect 14461 13475 14519 13481
rect 21652 13484 21916 13512
rect 13969 13447 14027 13453
rect 13969 13444 13981 13447
rect 13740 13416 13981 13444
rect 13969 13413 13981 13416
rect 14015 13444 14027 13447
rect 14185 13447 14243 13453
rect 14015 13413 14044 13444
rect 13969 13407 14044 13413
rect 14185 13413 14197 13447
rect 14231 13413 14243 13447
rect 14185 13407 14243 13413
rect 13357 13379 13415 13385
rect 13357 13345 13369 13379
rect 13403 13345 13415 13379
rect 13357 13339 13415 13345
rect 13541 13379 13599 13385
rect 13541 13345 13553 13379
rect 13587 13345 13599 13379
rect 14016 13376 14044 13407
rect 17494 13404 17500 13456
rect 17552 13404 17558 13456
rect 14277 13379 14335 13385
rect 14277 13376 14289 13379
rect 14016 13348 14289 13376
rect 13541 13339 13599 13345
rect 14277 13345 14289 13348
rect 14323 13345 14335 13379
rect 14277 13339 14335 13345
rect 14553 13379 14611 13385
rect 14553 13345 14565 13379
rect 14599 13345 14611 13379
rect 14553 13339 14611 13345
rect 10008 13212 10916 13240
rect 10008 13200 10014 13212
rect 12342 13200 12348 13252
rect 12400 13240 12406 13252
rect 13372 13240 13400 13339
rect 14568 13308 14596 13339
rect 17218 13336 17224 13388
rect 17276 13376 17282 13388
rect 17313 13379 17371 13385
rect 17313 13376 17325 13379
rect 17276 13348 17325 13376
rect 17276 13336 17282 13348
rect 17313 13345 17325 13348
rect 17359 13345 17371 13379
rect 17313 13339 17371 13345
rect 21450 13336 21456 13388
rect 21508 13336 21514 13388
rect 14016 13280 14596 13308
rect 14016 13240 14044 13280
rect 12400 13212 13400 13240
rect 13740 13212 14044 13240
rect 12400 13200 12406 13212
rect 2961 13175 3019 13181
rect 2961 13141 2973 13175
rect 3007 13172 3019 13175
rect 3418 13172 3424 13184
rect 3007 13144 3424 13172
rect 3007 13141 3019 13144
rect 2961 13135 3019 13141
rect 3418 13132 3424 13144
rect 3476 13132 3482 13184
rect 9674 13132 9680 13184
rect 9732 13132 9738 13184
rect 10410 13132 10416 13184
rect 10468 13132 10474 13184
rect 10502 13132 10508 13184
rect 10560 13132 10566 13184
rect 13354 13132 13360 13184
rect 13412 13172 13418 13184
rect 13740 13181 13768 13212
rect 13725 13175 13783 13181
rect 13725 13172 13737 13175
rect 13412 13144 13737 13172
rect 13412 13132 13418 13144
rect 13725 13141 13737 13144
rect 13771 13141 13783 13175
rect 13725 13135 13783 13141
rect 13814 13132 13820 13184
rect 13872 13132 13878 13184
rect 14016 13181 14044 13212
rect 17310 13200 17316 13252
rect 17368 13240 17374 13252
rect 19058 13240 19064 13252
rect 17368 13212 19064 13240
rect 17368 13200 17374 13212
rect 19058 13200 19064 13212
rect 19116 13200 19122 13252
rect 21652 13240 21680 13484
rect 21910 13472 21916 13484
rect 21968 13472 21974 13524
rect 21726 13404 21732 13456
rect 21784 13404 21790 13456
rect 22278 13404 22284 13456
rect 22336 13444 22342 13456
rect 22675 13447 22733 13453
rect 22675 13444 22687 13447
rect 22336 13416 22687 13444
rect 22336 13404 22342 13416
rect 22675 13413 22687 13416
rect 22721 13413 22733 13447
rect 22675 13407 22733 13413
rect 21744 13376 21772 13404
rect 21913 13379 21971 13385
rect 21744 13348 21864 13376
rect 21726 13268 21732 13320
rect 21784 13268 21790 13320
rect 21836 13308 21864 13348
rect 21913 13345 21925 13379
rect 21959 13376 21971 13379
rect 22189 13379 22247 13385
rect 22189 13376 22201 13379
rect 21959 13348 22201 13376
rect 21959 13345 21971 13348
rect 21913 13339 21971 13345
rect 22189 13345 22201 13348
rect 22235 13345 22247 13379
rect 22189 13339 22247 13345
rect 22373 13379 22431 13385
rect 22373 13345 22385 13379
rect 22419 13345 22431 13379
rect 22373 13339 22431 13345
rect 22388 13308 22416 13339
rect 22462 13336 22468 13388
rect 22520 13336 22526 13388
rect 22557 13379 22615 13385
rect 22557 13345 22569 13379
rect 22603 13345 22615 13379
rect 22557 13339 22615 13345
rect 21836 13280 22416 13308
rect 22097 13243 22155 13249
rect 22097 13240 22109 13243
rect 21652 13212 22109 13240
rect 22097 13209 22109 13212
rect 22143 13209 22155 13243
rect 22097 13203 22155 13209
rect 22186 13200 22192 13252
rect 22244 13240 22250 13252
rect 22572 13240 22600 13339
rect 22830 13268 22836 13320
rect 22888 13268 22894 13320
rect 22244 13212 22600 13240
rect 22244 13200 22250 13212
rect 14001 13175 14059 13181
rect 14001 13141 14013 13175
rect 14047 13141 14059 13175
rect 14001 13135 14059 13141
rect 14274 13132 14280 13184
rect 14332 13132 14338 13184
rect 17681 13175 17739 13181
rect 17681 13141 17693 13175
rect 17727 13172 17739 13175
rect 17770 13172 17776 13184
rect 17727 13144 17776 13172
rect 17727 13141 17739 13144
rect 17681 13135 17739 13141
rect 17770 13132 17776 13144
rect 17828 13132 17834 13184
rect 21913 13175 21971 13181
rect 21913 13141 21925 13175
rect 21959 13172 21971 13175
rect 22002 13172 22008 13184
rect 21959 13144 22008 13172
rect 21959 13141 21971 13144
rect 21913 13135 21971 13141
rect 22002 13132 22008 13144
rect 22060 13132 22066 13184
rect 552 13082 23368 13104
rect 552 13030 3662 13082
rect 3714 13030 3726 13082
rect 3778 13030 3790 13082
rect 3842 13030 3854 13082
rect 3906 13030 3918 13082
rect 3970 13030 23368 13082
rect 552 13008 23368 13030
rect 8754 12928 8760 12980
rect 8812 12968 8818 12980
rect 9398 12968 9404 12980
rect 8812 12940 9404 12968
rect 8812 12928 8818 12940
rect 9398 12928 9404 12940
rect 9456 12928 9462 12980
rect 12434 12968 12440 12980
rect 12084 12940 12440 12968
rect 9125 12903 9183 12909
rect 6932 12872 7420 12900
rect 6932 12844 6960 12872
rect 5169 12835 5227 12841
rect 5169 12801 5181 12835
rect 5215 12832 5227 12835
rect 5258 12832 5264 12844
rect 5215 12804 5264 12832
rect 5215 12801 5227 12804
rect 5169 12795 5227 12801
rect 5258 12792 5264 12804
rect 5316 12792 5322 12844
rect 6914 12792 6920 12844
rect 6972 12792 6978 12844
rect 7190 12792 7196 12844
rect 7248 12792 7254 12844
rect 4893 12767 4951 12773
rect 4893 12733 4905 12767
rect 4939 12764 4951 12767
rect 4982 12764 4988 12776
rect 4939 12736 4988 12764
rect 4939 12733 4951 12736
rect 4893 12727 4951 12733
rect 4982 12724 4988 12736
rect 5040 12764 5046 12776
rect 5350 12764 5356 12776
rect 5040 12736 5356 12764
rect 5040 12724 5046 12736
rect 5350 12724 5356 12736
rect 5408 12724 5414 12776
rect 7392 12773 7420 12872
rect 9125 12869 9137 12903
rect 9171 12900 9183 12903
rect 9674 12900 9680 12912
rect 9171 12872 9680 12900
rect 9171 12869 9183 12872
rect 9125 12863 9183 12869
rect 9674 12860 9680 12872
rect 9732 12860 9738 12912
rect 8570 12792 8576 12844
rect 8628 12832 8634 12844
rect 8757 12835 8815 12841
rect 8757 12832 8769 12835
rect 8628 12804 8769 12832
rect 8628 12792 8634 12804
rect 8757 12801 8769 12804
rect 8803 12801 8815 12835
rect 8757 12795 8815 12801
rect 8864 12804 9260 12832
rect 8864 12776 8892 12804
rect 6825 12767 6883 12773
rect 6825 12733 6837 12767
rect 6871 12764 6883 12767
rect 7285 12767 7343 12773
rect 7285 12764 7297 12767
rect 6871 12736 7297 12764
rect 6871 12733 6883 12736
rect 6825 12727 6883 12733
rect 7285 12733 7297 12736
rect 7331 12733 7343 12767
rect 7285 12727 7343 12733
rect 7378 12767 7436 12773
rect 7378 12733 7390 12767
rect 7424 12733 7436 12767
rect 7378 12727 7436 12733
rect 8481 12767 8539 12773
rect 8481 12733 8493 12767
rect 8527 12764 8539 12767
rect 8662 12764 8668 12776
rect 8527 12736 8668 12764
rect 8527 12733 8539 12736
rect 8481 12727 8539 12733
rect 7300 12696 7328 12727
rect 8662 12724 8668 12736
rect 8720 12764 8726 12776
rect 8846 12764 8852 12776
rect 8720 12736 8852 12764
rect 8720 12724 8726 12736
rect 8846 12724 8852 12736
rect 8904 12724 8910 12776
rect 9232 12773 9260 12804
rect 10410 12792 10416 12844
rect 10468 12832 10474 12844
rect 12084 12841 12112 12940
rect 12434 12928 12440 12940
rect 12492 12928 12498 12980
rect 12526 12928 12532 12980
rect 12584 12968 12590 12980
rect 12805 12971 12863 12977
rect 12805 12968 12817 12971
rect 12584 12940 12817 12968
rect 12584 12928 12590 12940
rect 12805 12937 12817 12940
rect 12851 12968 12863 12971
rect 13262 12968 13268 12980
rect 12851 12940 13268 12968
rect 12851 12937 12863 12940
rect 12805 12931 12863 12937
rect 13262 12928 13268 12940
rect 13320 12928 13326 12980
rect 13725 12971 13783 12977
rect 13725 12937 13737 12971
rect 13771 12968 13783 12971
rect 14274 12968 14280 12980
rect 13771 12940 14280 12968
rect 13771 12937 13783 12940
rect 13725 12931 13783 12937
rect 14274 12928 14280 12940
rect 14332 12928 14338 12980
rect 17681 12971 17739 12977
rect 17681 12937 17693 12971
rect 17727 12968 17739 12971
rect 17770 12968 17776 12980
rect 17727 12940 17776 12968
rect 17727 12937 17739 12940
rect 17681 12931 17739 12937
rect 17770 12928 17776 12940
rect 17828 12928 17834 12980
rect 18233 12971 18291 12977
rect 18233 12937 18245 12971
rect 18279 12968 18291 12971
rect 18322 12968 18328 12980
rect 18279 12940 18328 12968
rect 18279 12937 18291 12940
rect 18233 12931 18291 12937
rect 18322 12928 18328 12940
rect 18380 12928 18386 12980
rect 18417 12971 18475 12977
rect 18417 12937 18429 12971
rect 18463 12968 18475 12971
rect 20162 12968 20168 12980
rect 18463 12940 20168 12968
rect 18463 12937 18475 12940
rect 18417 12931 18475 12937
rect 20162 12928 20168 12940
rect 20220 12928 20226 12980
rect 21726 12928 21732 12980
rect 21784 12928 21790 12980
rect 19518 12900 19524 12912
rect 12728 12872 19524 12900
rect 12069 12835 12127 12841
rect 12069 12832 12081 12835
rect 10468 12804 12081 12832
rect 10468 12792 10474 12804
rect 12069 12801 12081 12804
rect 12115 12801 12127 12835
rect 12069 12795 12127 12801
rect 12161 12835 12219 12841
rect 12161 12801 12173 12835
rect 12207 12832 12219 12835
rect 12250 12832 12256 12844
rect 12207 12804 12256 12832
rect 12207 12801 12219 12804
rect 12161 12795 12219 12801
rect 12250 12792 12256 12804
rect 12308 12832 12314 12844
rect 12728 12832 12756 12872
rect 19518 12860 19524 12872
rect 19576 12860 19582 12912
rect 21634 12860 21640 12912
rect 21692 12900 21698 12912
rect 21692 12872 22048 12900
rect 21692 12860 21698 12872
rect 12308 12804 12756 12832
rect 12308 12792 12314 12804
rect 12802 12792 12808 12844
rect 12860 12832 12866 12844
rect 12860 12804 13032 12832
rect 12860 12792 12866 12804
rect 8941 12767 8999 12773
rect 8941 12733 8953 12767
rect 8987 12733 8999 12767
rect 8941 12727 8999 12733
rect 9217 12767 9275 12773
rect 9217 12733 9229 12767
rect 9263 12733 9275 12767
rect 9217 12727 9275 12733
rect 8386 12696 8392 12708
rect 7300 12668 8392 12696
rect 8386 12656 8392 12668
rect 8444 12656 8450 12708
rect 4246 12588 4252 12640
rect 4304 12628 4310 12640
rect 4525 12631 4583 12637
rect 4525 12628 4537 12631
rect 4304 12600 4537 12628
rect 4304 12588 4310 12600
rect 4525 12597 4537 12600
rect 4571 12597 4583 12631
rect 4525 12591 4583 12597
rect 4798 12588 4804 12640
rect 4856 12628 4862 12640
rect 4985 12631 5043 12637
rect 4985 12628 4997 12631
rect 4856 12600 4997 12628
rect 4856 12588 4862 12600
rect 4985 12597 4997 12600
rect 5031 12597 5043 12631
rect 4985 12591 5043 12597
rect 7653 12631 7711 12637
rect 7653 12597 7665 12631
rect 7699 12628 7711 12631
rect 7926 12628 7932 12640
rect 7699 12600 7932 12628
rect 7699 12597 7711 12600
rect 7653 12591 7711 12597
rect 7926 12588 7932 12600
rect 7984 12628 7990 12640
rect 8956 12628 8984 12727
rect 9398 12724 9404 12776
rect 9456 12724 9462 12776
rect 11882 12724 11888 12776
rect 11940 12724 11946 12776
rect 11977 12767 12035 12773
rect 11977 12733 11989 12767
rect 12023 12764 12035 12767
rect 12345 12767 12403 12773
rect 12345 12764 12357 12767
rect 12023 12736 12357 12764
rect 12023 12733 12035 12736
rect 11977 12727 12035 12733
rect 12345 12733 12357 12736
rect 12391 12733 12403 12767
rect 12345 12727 12403 12733
rect 10686 12656 10692 12708
rect 10744 12696 10750 12708
rect 11992 12696 12020 12727
rect 12434 12724 12440 12776
rect 12492 12724 12498 12776
rect 12621 12767 12679 12773
rect 12621 12733 12633 12767
rect 12667 12764 12679 12767
rect 12710 12764 12716 12776
rect 12667 12736 12716 12764
rect 12667 12733 12679 12736
rect 12621 12727 12679 12733
rect 12636 12696 12664 12727
rect 12710 12724 12716 12736
rect 12768 12724 12774 12776
rect 13004 12773 13032 12804
rect 13446 12792 13452 12844
rect 13504 12832 13510 12844
rect 13541 12835 13599 12841
rect 13541 12832 13553 12835
rect 13504 12804 13553 12832
rect 13504 12792 13510 12804
rect 13541 12801 13553 12804
rect 13587 12832 13599 12835
rect 13587 12804 15240 12832
rect 13587 12801 13599 12804
rect 13541 12795 13599 12801
rect 12897 12767 12955 12773
rect 12897 12733 12909 12767
rect 12943 12733 12955 12767
rect 12897 12727 12955 12733
rect 12990 12767 13048 12773
rect 12990 12733 13002 12767
rect 13036 12733 13048 12767
rect 12990 12727 13048 12733
rect 12912 12696 12940 12727
rect 13814 12724 13820 12776
rect 13872 12724 13878 12776
rect 15212 12764 15240 12804
rect 15286 12792 15292 12844
rect 15344 12832 15350 12844
rect 15381 12835 15439 12841
rect 15381 12832 15393 12835
rect 15344 12804 15393 12832
rect 15344 12792 15350 12804
rect 15381 12801 15393 12804
rect 15427 12801 15439 12835
rect 15381 12795 15439 12801
rect 15473 12835 15531 12841
rect 15473 12801 15485 12835
rect 15519 12832 15531 12835
rect 17310 12832 17316 12844
rect 15519 12804 17316 12832
rect 15519 12801 15531 12804
rect 15473 12795 15531 12801
rect 15488 12764 15516 12795
rect 17310 12792 17316 12804
rect 17368 12792 17374 12844
rect 17494 12832 17500 12844
rect 17420 12804 17500 12832
rect 15212 12736 15516 12764
rect 17218 12724 17224 12776
rect 17276 12724 17282 12776
rect 17420 12773 17448 12804
rect 17494 12792 17500 12804
rect 17552 12792 17558 12844
rect 18046 12792 18052 12844
rect 18104 12792 18110 12844
rect 21818 12792 21824 12844
rect 21876 12832 21882 12844
rect 21876 12804 21956 12832
rect 21876 12792 21882 12804
rect 17405 12767 17463 12773
rect 17405 12733 17417 12767
rect 17451 12733 17463 12767
rect 18138 12764 18144 12776
rect 17405 12727 17463 12733
rect 17512 12736 18144 12764
rect 10744 12668 12020 12696
rect 12084 12668 12664 12696
rect 12728 12668 12940 12696
rect 15289 12699 15347 12705
rect 10744 12656 10750 12668
rect 7984 12600 8984 12628
rect 7984 12588 7990 12600
rect 9398 12588 9404 12640
rect 9456 12588 9462 12640
rect 11698 12588 11704 12640
rect 11756 12588 11762 12640
rect 11882 12588 11888 12640
rect 11940 12628 11946 12640
rect 12084 12628 12112 12668
rect 11940 12600 12112 12628
rect 11940 12588 11946 12600
rect 12434 12588 12440 12640
rect 12492 12628 12498 12640
rect 12728 12628 12756 12668
rect 15289 12665 15301 12699
rect 15335 12696 15347 12699
rect 15930 12696 15936 12708
rect 15335 12668 15936 12696
rect 15335 12665 15347 12668
rect 15289 12659 15347 12665
rect 15930 12656 15936 12668
rect 15988 12656 15994 12708
rect 17512 12705 17540 12736
rect 18138 12724 18144 12736
rect 18196 12724 18202 12776
rect 18230 12724 18236 12776
rect 18288 12724 18294 12776
rect 17497 12699 17555 12705
rect 17497 12665 17509 12699
rect 17543 12665 17555 12699
rect 17497 12659 17555 12665
rect 17954 12656 17960 12708
rect 18012 12656 18018 12708
rect 21928 12705 21956 12804
rect 22020 12773 22048 12872
rect 22005 12767 22063 12773
rect 22005 12733 22017 12767
rect 22051 12733 22063 12767
rect 22005 12727 22063 12733
rect 21729 12699 21787 12705
rect 21729 12665 21741 12699
rect 21775 12665 21787 12699
rect 21729 12659 21787 12665
rect 21913 12699 21971 12705
rect 21913 12665 21925 12699
rect 21959 12696 21971 12699
rect 22462 12696 22468 12708
rect 21959 12668 22468 12696
rect 21959 12665 21971 12668
rect 21913 12659 21971 12665
rect 12492 12600 12756 12628
rect 12492 12588 12498 12600
rect 13262 12588 13268 12640
rect 13320 12588 13326 12640
rect 13541 12631 13599 12637
rect 13541 12597 13553 12631
rect 13587 12628 13599 12631
rect 14366 12628 14372 12640
rect 13587 12600 14372 12628
rect 13587 12597 13599 12600
rect 13541 12591 13599 12597
rect 14366 12588 14372 12600
rect 14424 12588 14430 12640
rect 14918 12588 14924 12640
rect 14976 12588 14982 12640
rect 17405 12631 17463 12637
rect 17405 12597 17417 12631
rect 17451 12628 17463 12631
rect 17678 12628 17684 12640
rect 17736 12637 17742 12640
rect 17736 12631 17755 12637
rect 17451 12600 17684 12628
rect 17451 12597 17463 12600
rect 17405 12591 17463 12597
rect 17678 12588 17684 12600
rect 17743 12597 17755 12631
rect 17736 12591 17755 12597
rect 17865 12631 17923 12637
rect 17865 12597 17877 12631
rect 17911 12628 17923 12631
rect 18874 12628 18880 12640
rect 17911 12600 18880 12628
rect 17911 12597 17923 12600
rect 17865 12591 17923 12597
rect 17736 12588 17742 12591
rect 18874 12588 18880 12600
rect 18932 12588 18938 12640
rect 21744 12628 21772 12659
rect 22462 12656 22468 12668
rect 22520 12656 22526 12708
rect 22186 12628 22192 12640
rect 21744 12600 22192 12628
rect 22186 12588 22192 12600
rect 22244 12588 22250 12640
rect 552 12538 23368 12560
rect 552 12486 4322 12538
rect 4374 12486 4386 12538
rect 4438 12486 4450 12538
rect 4502 12486 4514 12538
rect 4566 12486 4578 12538
rect 4630 12486 23368 12538
rect 552 12464 23368 12486
rect 2774 12384 2780 12436
rect 2832 12424 2838 12436
rect 3421 12427 3479 12433
rect 3421 12424 3433 12427
rect 2832 12396 3433 12424
rect 2832 12384 2838 12396
rect 3421 12393 3433 12396
rect 3467 12393 3479 12427
rect 3421 12387 3479 12393
rect 5350 12384 5356 12436
rect 5408 12384 5414 12436
rect 9398 12384 9404 12436
rect 9456 12424 9462 12436
rect 10337 12427 10395 12433
rect 9456 12396 10180 12424
rect 9456 12384 9462 12396
rect 4246 12365 4252 12368
rect 4240 12356 4252 12365
rect 4207 12328 4252 12356
rect 4240 12319 4252 12328
rect 4246 12316 4252 12319
rect 4304 12316 4310 12368
rect 8570 12316 8576 12368
rect 8628 12356 8634 12368
rect 8665 12359 8723 12365
rect 8665 12356 8677 12359
rect 8628 12328 8677 12356
rect 8628 12316 8634 12328
rect 8665 12325 8677 12328
rect 8711 12325 8723 12359
rect 8665 12319 8723 12325
rect 8846 12316 8852 12368
rect 8904 12316 8910 12368
rect 9674 12316 9680 12368
rect 9732 12316 9738 12368
rect 9784 12365 9812 12396
rect 10152 12365 10180 12396
rect 10337 12393 10349 12427
rect 10383 12424 10395 12427
rect 10383 12396 10640 12424
rect 10383 12393 10395 12396
rect 10337 12387 10395 12393
rect 9769 12359 9827 12365
rect 9769 12325 9781 12359
rect 9815 12325 9827 12359
rect 9769 12319 9827 12325
rect 10137 12359 10195 12365
rect 10137 12325 10149 12359
rect 10183 12325 10195 12359
rect 10137 12319 10195 12325
rect 3973 12291 4031 12297
rect 3973 12257 3985 12291
rect 4019 12288 4031 12291
rect 4614 12288 4620 12300
rect 4019 12260 4620 12288
rect 4019 12257 4031 12260
rect 3973 12251 4031 12257
rect 4614 12248 4620 12260
rect 4672 12248 4678 12300
rect 7190 12248 7196 12300
rect 7248 12288 7254 12300
rect 7285 12291 7343 12297
rect 7285 12288 7297 12291
rect 7248 12260 7297 12288
rect 7248 12248 7254 12260
rect 7285 12257 7297 12260
rect 7331 12257 7343 12291
rect 7285 12251 7343 12257
rect 7374 12248 7380 12300
rect 7432 12288 7438 12300
rect 7469 12291 7527 12297
rect 7469 12288 7481 12291
rect 7432 12260 7481 12288
rect 7432 12248 7438 12260
rect 7469 12257 7481 12260
rect 7515 12257 7527 12291
rect 7469 12251 7527 12257
rect 8021 12291 8079 12297
rect 8021 12257 8033 12291
rect 8067 12257 8079 12291
rect 8021 12251 8079 12257
rect 3234 12180 3240 12232
rect 3292 12180 3298 12232
rect 3326 12180 3332 12232
rect 3384 12180 3390 12232
rect 7834 12220 7840 12232
rect 7484 12192 7840 12220
rect 7484 12161 7512 12192
rect 7834 12180 7840 12192
rect 7892 12220 7898 12232
rect 8036 12220 8064 12251
rect 8202 12248 8208 12300
rect 8260 12248 8266 12300
rect 8481 12291 8539 12297
rect 8481 12257 8493 12291
rect 8527 12288 8539 12291
rect 8754 12288 8760 12300
rect 8527 12260 8760 12288
rect 8527 12257 8539 12260
rect 8481 12251 8539 12257
rect 8754 12248 8760 12260
rect 8812 12288 8818 12300
rect 9033 12291 9091 12297
rect 9033 12288 9045 12291
rect 8812 12260 9045 12288
rect 8812 12248 8818 12260
rect 9033 12257 9045 12260
rect 9079 12257 9091 12291
rect 9033 12251 9091 12257
rect 9585 12291 9643 12297
rect 9585 12257 9597 12291
rect 9631 12257 9643 12291
rect 9585 12251 9643 12257
rect 7892 12192 8064 12220
rect 8113 12223 8171 12229
rect 7892 12180 7898 12192
rect 8113 12189 8125 12223
rect 8159 12220 8171 12223
rect 9600 12220 9628 12251
rect 9950 12248 9956 12300
rect 10008 12248 10014 12300
rect 10045 12291 10103 12297
rect 10045 12257 10057 12291
rect 10091 12288 10103 12291
rect 10226 12288 10232 12300
rect 10091 12260 10232 12288
rect 10091 12257 10103 12260
rect 10045 12251 10103 12257
rect 10226 12248 10232 12260
rect 10284 12288 10290 12300
rect 10502 12288 10508 12300
rect 10284 12260 10508 12288
rect 10284 12248 10290 12260
rect 10502 12248 10508 12260
rect 10560 12248 10566 12300
rect 10612 12220 10640 12396
rect 12434 12384 12440 12436
rect 12492 12384 12498 12436
rect 16684 12396 17448 12424
rect 16684 12368 16712 12396
rect 14820 12359 14878 12365
rect 14820 12325 14832 12359
rect 14866 12356 14878 12359
rect 14918 12356 14924 12368
rect 14866 12328 14924 12356
rect 14866 12325 14878 12328
rect 14820 12319 14878 12325
rect 14918 12316 14924 12328
rect 14976 12316 14982 12368
rect 16666 12316 16672 12368
rect 16724 12316 16730 12368
rect 17420 12365 17448 12396
rect 17770 12384 17776 12436
rect 17828 12384 17834 12436
rect 18049 12427 18107 12433
rect 18049 12393 18061 12427
rect 18095 12424 18107 12427
rect 18230 12424 18236 12436
rect 18095 12396 18236 12424
rect 18095 12393 18107 12396
rect 18049 12387 18107 12393
rect 18230 12384 18236 12396
rect 18288 12384 18294 12436
rect 18322 12384 18328 12436
rect 18380 12424 18386 12436
rect 19061 12427 19119 12433
rect 19061 12424 19073 12427
rect 18380 12396 19073 12424
rect 18380 12384 18386 12396
rect 19061 12393 19073 12396
rect 19107 12393 19119 12427
rect 19061 12387 19119 12393
rect 22738 12384 22744 12436
rect 22796 12424 22802 12436
rect 22833 12427 22891 12433
rect 22833 12424 22845 12427
rect 22796 12396 22845 12424
rect 22796 12384 22802 12396
rect 22833 12393 22845 12396
rect 22879 12393 22891 12427
rect 22833 12387 22891 12393
rect 16885 12359 16943 12365
rect 16885 12325 16897 12359
rect 16931 12356 16943 12359
rect 17405 12359 17463 12365
rect 16931 12328 17172 12356
rect 16931 12325 16943 12328
rect 16885 12319 16943 12325
rect 17144 12300 17172 12328
rect 17405 12325 17417 12359
rect 17451 12325 17463 12359
rect 17405 12319 17463 12325
rect 17957 12359 18015 12365
rect 17957 12325 17969 12359
rect 18003 12356 18015 12359
rect 18138 12356 18144 12368
rect 18003 12328 18144 12356
rect 18003 12325 18015 12328
rect 17957 12319 18015 12325
rect 18138 12316 18144 12328
rect 18196 12316 18202 12368
rect 18874 12316 18880 12368
rect 18932 12316 18938 12368
rect 20257 12359 20315 12365
rect 20257 12325 20269 12359
rect 20303 12325 20315 12359
rect 20257 12319 20315 12325
rect 12342 12248 12348 12300
rect 12400 12248 12406 12300
rect 12526 12248 12532 12300
rect 12584 12248 12590 12300
rect 13262 12248 13268 12300
rect 13320 12248 13326 12300
rect 13354 12248 13360 12300
rect 13412 12248 13418 12300
rect 13446 12248 13452 12300
rect 13504 12288 13510 12300
rect 14274 12288 14280 12300
rect 13504 12260 14280 12288
rect 13504 12248 13510 12260
rect 14274 12248 14280 12260
rect 14332 12248 14338 12300
rect 17126 12248 17132 12300
rect 17184 12248 17190 12300
rect 17218 12248 17224 12300
rect 17276 12248 17282 12300
rect 17678 12248 17684 12300
rect 17736 12248 17742 12300
rect 18414 12248 18420 12300
rect 18472 12248 18478 12300
rect 18693 12291 18751 12297
rect 18693 12288 18705 12291
rect 18616 12260 18705 12288
rect 8159 12192 10640 12220
rect 8159 12189 8171 12192
rect 8113 12183 8171 12189
rect 13538 12180 13544 12232
rect 13596 12180 13602 12232
rect 14550 12180 14556 12232
rect 14608 12180 14614 12232
rect 7469 12155 7527 12161
rect 7469 12121 7481 12155
rect 7515 12121 7527 12155
rect 7469 12115 7527 12121
rect 9401 12155 9459 12161
rect 9401 12121 9413 12155
rect 9447 12152 9459 12155
rect 10686 12152 10692 12164
rect 9447 12124 10692 12152
rect 9447 12121 9459 12124
rect 9401 12115 9459 12121
rect 10686 12112 10692 12124
rect 10744 12112 10750 12164
rect 3789 12087 3847 12093
rect 3789 12053 3801 12087
rect 3835 12084 3847 12087
rect 4338 12084 4344 12096
rect 3835 12056 4344 12084
rect 3835 12053 3847 12056
rect 3789 12047 3847 12053
rect 4338 12044 4344 12056
rect 4396 12044 4402 12096
rect 8297 12087 8355 12093
rect 8297 12053 8309 12087
rect 8343 12084 8355 12087
rect 8386 12084 8392 12096
rect 8343 12056 8392 12084
rect 8343 12053 8355 12056
rect 8297 12047 8355 12053
rect 8386 12044 8392 12056
rect 8444 12044 8450 12096
rect 9217 12087 9275 12093
rect 9217 12053 9229 12087
rect 9263 12084 9275 12087
rect 9306 12084 9312 12096
rect 9263 12056 9312 12084
rect 9263 12053 9275 12056
rect 9217 12047 9275 12053
rect 9306 12044 9312 12056
rect 9364 12044 9370 12096
rect 9674 12044 9680 12096
rect 9732 12084 9738 12096
rect 10321 12087 10379 12093
rect 10321 12084 10333 12087
rect 9732 12056 10333 12084
rect 9732 12044 9738 12056
rect 10321 12053 10333 12056
rect 10367 12053 10379 12087
rect 10321 12047 10379 12053
rect 10502 12044 10508 12096
rect 10560 12044 10566 12096
rect 13078 12044 13084 12096
rect 13136 12044 13142 12096
rect 14568 12084 14596 12180
rect 17236 12152 17264 12248
rect 18506 12180 18512 12232
rect 18564 12180 18570 12232
rect 16868 12124 17264 12152
rect 17957 12155 18015 12161
rect 14918 12084 14924 12096
rect 14568 12056 14924 12084
rect 14918 12044 14924 12056
rect 14976 12044 14982 12096
rect 15930 12044 15936 12096
rect 15988 12084 15994 12096
rect 16114 12084 16120 12096
rect 15988 12056 16120 12084
rect 15988 12044 15994 12056
rect 16114 12044 16120 12056
rect 16172 12044 16178 12096
rect 16574 12044 16580 12096
rect 16632 12084 16638 12096
rect 16868 12093 16896 12124
rect 17957 12121 17969 12155
rect 18003 12152 18015 12155
rect 18616 12152 18644 12260
rect 18693 12257 18705 12260
rect 18739 12257 18751 12291
rect 20272 12288 20300 12319
rect 20346 12316 20352 12368
rect 20404 12356 20410 12368
rect 20457 12359 20515 12365
rect 20457 12356 20469 12359
rect 20404 12328 20469 12356
rect 20404 12316 20410 12328
rect 20457 12325 20469 12328
rect 20503 12325 20515 12359
rect 22756 12356 22784 12384
rect 20457 12319 20515 12325
rect 21744 12328 22784 12356
rect 20717 12291 20775 12297
rect 20717 12288 20729 12291
rect 20272 12260 20729 12288
rect 18693 12251 18751 12257
rect 20717 12257 20729 12260
rect 20763 12257 20775 12291
rect 20717 12251 20775 12257
rect 20901 12291 20959 12297
rect 20901 12257 20913 12291
rect 20947 12288 20959 12291
rect 21542 12288 21548 12300
rect 20947 12260 21548 12288
rect 20947 12257 20959 12260
rect 20901 12251 20959 12257
rect 20732 12220 20760 12251
rect 21542 12248 21548 12260
rect 21600 12248 21606 12300
rect 21744 12297 21772 12328
rect 21729 12291 21787 12297
rect 21729 12257 21741 12291
rect 21775 12257 21787 12291
rect 21729 12251 21787 12257
rect 21821 12291 21879 12297
rect 21821 12257 21833 12291
rect 21867 12288 21879 12291
rect 21910 12288 21916 12300
rect 21867 12260 21916 12288
rect 21867 12257 21879 12260
rect 21821 12251 21879 12257
rect 21910 12248 21916 12260
rect 21968 12248 21974 12300
rect 22094 12248 22100 12300
rect 22152 12288 22158 12300
rect 22281 12291 22339 12297
rect 22281 12288 22293 12291
rect 22152 12260 22293 12288
rect 22152 12248 22158 12260
rect 22281 12257 22293 12260
rect 22327 12257 22339 12291
rect 22281 12251 22339 12257
rect 23014 12248 23020 12300
rect 23072 12248 23078 12300
rect 20990 12220 20996 12232
rect 20732 12192 20996 12220
rect 20990 12180 20996 12192
rect 21048 12180 21054 12232
rect 18003 12124 18644 12152
rect 18003 12121 18015 12124
rect 17957 12115 18015 12121
rect 21542 12112 21548 12164
rect 21600 12152 21606 12164
rect 22097 12155 22155 12161
rect 22097 12152 22109 12155
rect 21600 12124 22109 12152
rect 21600 12112 21606 12124
rect 22097 12121 22109 12124
rect 22143 12121 22155 12155
rect 22097 12115 22155 12121
rect 16853 12087 16911 12093
rect 16853 12084 16865 12087
rect 16632 12056 16865 12084
rect 16632 12044 16638 12056
rect 16853 12053 16865 12056
rect 16899 12053 16911 12087
rect 16853 12047 16911 12053
rect 17034 12044 17040 12096
rect 17092 12044 17098 12096
rect 17310 12044 17316 12096
rect 17368 12084 17374 12096
rect 17405 12087 17463 12093
rect 17405 12084 17417 12087
rect 17368 12056 17417 12084
rect 17368 12044 17374 12056
rect 17405 12053 17417 12056
rect 17451 12053 17463 12087
rect 17405 12047 17463 12053
rect 19518 12044 19524 12096
rect 19576 12084 19582 12096
rect 20441 12087 20499 12093
rect 20441 12084 20453 12087
rect 19576 12056 20453 12084
rect 19576 12044 19582 12056
rect 20441 12053 20453 12056
rect 20487 12053 20499 12087
rect 20441 12047 20499 12053
rect 20625 12087 20683 12093
rect 20625 12053 20637 12087
rect 20671 12084 20683 12087
rect 20714 12084 20720 12096
rect 20671 12056 20720 12084
rect 20671 12053 20683 12056
rect 20625 12047 20683 12053
rect 20714 12044 20720 12056
rect 20772 12044 20778 12096
rect 22002 12044 22008 12096
rect 22060 12044 22066 12096
rect 552 11994 23368 12016
rect 552 11942 3662 11994
rect 3714 11942 3726 11994
rect 3778 11942 3790 11994
rect 3842 11942 3854 11994
rect 3906 11942 3918 11994
rect 3970 11942 23368 11994
rect 552 11920 23368 11942
rect 3237 11883 3295 11889
rect 3237 11849 3249 11883
rect 3283 11880 3295 11883
rect 3326 11880 3332 11892
rect 3283 11852 3332 11880
rect 3283 11849 3295 11852
rect 3237 11843 3295 11849
rect 3326 11840 3332 11852
rect 3384 11840 3390 11892
rect 10137 11883 10195 11889
rect 10137 11849 10149 11883
rect 10183 11880 10195 11883
rect 10226 11880 10232 11892
rect 10183 11852 10232 11880
rect 10183 11849 10195 11852
rect 10137 11843 10195 11849
rect 10226 11840 10232 11852
rect 10284 11840 10290 11892
rect 16206 11840 16212 11892
rect 16264 11840 16270 11892
rect 16393 11883 16451 11889
rect 16393 11849 16405 11883
rect 16439 11880 16451 11883
rect 16574 11880 16580 11892
rect 16439 11852 16580 11880
rect 16439 11849 16451 11852
rect 16393 11843 16451 11849
rect 16574 11840 16580 11852
rect 16632 11840 16638 11892
rect 16669 11883 16727 11889
rect 16669 11849 16681 11883
rect 16715 11880 16727 11883
rect 17126 11880 17132 11892
rect 16715 11852 17132 11880
rect 16715 11849 16727 11852
rect 16669 11843 16727 11849
rect 17126 11840 17132 11852
rect 17184 11840 17190 11892
rect 17681 11883 17739 11889
rect 17681 11849 17693 11883
rect 17727 11880 17739 11883
rect 18046 11880 18052 11892
rect 17727 11852 18052 11880
rect 17727 11849 17739 11852
rect 17681 11843 17739 11849
rect 18046 11840 18052 11852
rect 18104 11840 18110 11892
rect 19518 11840 19524 11892
rect 19576 11840 19582 11892
rect 20073 11883 20131 11889
rect 20073 11849 20085 11883
rect 20119 11880 20131 11883
rect 20346 11880 20352 11892
rect 20119 11852 20352 11880
rect 20119 11849 20131 11852
rect 20073 11843 20131 11849
rect 20346 11840 20352 11852
rect 20404 11840 20410 11892
rect 20806 11880 20812 11892
rect 20456 11852 20812 11880
rect 7009 11815 7067 11821
rect 4816 11784 6914 11812
rect 4614 11704 4620 11756
rect 4672 11744 4678 11756
rect 4816 11744 4844 11784
rect 4672 11716 4844 11744
rect 4672 11704 4678 11716
rect 4890 11704 4896 11756
rect 4948 11744 4954 11756
rect 5169 11747 5227 11753
rect 5169 11744 5181 11747
rect 4948 11716 5181 11744
rect 4948 11704 4954 11716
rect 5169 11713 5181 11716
rect 5215 11713 5227 11747
rect 5169 11707 5227 11713
rect 5258 11704 5264 11756
rect 5316 11704 5322 11756
rect 6886 11744 6914 11784
rect 7009 11781 7021 11815
rect 7055 11812 7067 11815
rect 7558 11812 7564 11824
rect 7055 11784 7564 11812
rect 7055 11781 7067 11784
rect 7009 11775 7067 11781
rect 7558 11772 7564 11784
rect 7616 11772 7622 11824
rect 9858 11744 9864 11756
rect 6886 11716 9864 11744
rect 9858 11704 9864 11716
rect 9916 11704 9922 11756
rect 10321 11747 10379 11753
rect 10321 11713 10333 11747
rect 10367 11744 10379 11747
rect 10502 11744 10508 11756
rect 10367 11716 10508 11744
rect 10367 11713 10379 11716
rect 10321 11707 10379 11713
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 10686 11704 10692 11756
rect 10744 11704 10750 11756
rect 14918 11704 14924 11756
rect 14976 11704 14982 11756
rect 16224 11744 16252 11840
rect 20165 11815 20223 11821
rect 20165 11781 20177 11815
rect 20211 11812 20223 11815
rect 20456 11812 20484 11852
rect 20806 11840 20812 11852
rect 20864 11840 20870 11892
rect 21174 11840 21180 11892
rect 21232 11880 21238 11892
rect 21232 11852 21588 11880
rect 21232 11840 21238 11852
rect 20211 11784 20484 11812
rect 20211 11781 20223 11784
rect 20165 11775 20223 11781
rect 16761 11747 16819 11753
rect 16761 11744 16773 11747
rect 16224 11716 16773 11744
rect 16761 11713 16773 11716
rect 16807 11713 16819 11747
rect 16761 11707 16819 11713
rect 17034 11704 17040 11756
rect 17092 11744 17098 11756
rect 17092 11716 17540 11744
rect 17092 11704 17098 11716
rect 4338 11636 4344 11688
rect 4396 11685 4402 11688
rect 4396 11676 4408 11685
rect 4396 11648 4441 11676
rect 4396 11639 4408 11648
rect 4396 11636 4402 11639
rect 7190 11636 7196 11688
rect 7248 11636 7254 11688
rect 7285 11679 7343 11685
rect 7285 11645 7297 11679
rect 7331 11676 7343 11679
rect 7374 11676 7380 11688
rect 7331 11648 7380 11676
rect 7331 11645 7343 11648
rect 7285 11639 7343 11645
rect 7374 11636 7380 11648
rect 7432 11636 7438 11688
rect 7926 11636 7932 11688
rect 7984 11636 7990 11688
rect 8113 11679 8171 11685
rect 8113 11645 8125 11679
rect 8159 11676 8171 11679
rect 8386 11676 8392 11688
rect 8159 11648 8392 11676
rect 8159 11645 8171 11648
rect 8113 11639 8171 11645
rect 8386 11636 8392 11648
rect 8444 11636 8450 11688
rect 9306 11636 9312 11688
rect 9364 11636 9370 11688
rect 9398 11636 9404 11688
rect 9456 11636 9462 11688
rect 9950 11636 9956 11688
rect 10008 11676 10014 11688
rect 10045 11679 10103 11685
rect 10045 11676 10057 11679
rect 10008 11648 10057 11676
rect 10008 11636 10014 11648
rect 10045 11645 10057 11648
rect 10091 11645 10103 11679
rect 10045 11639 10103 11645
rect 10597 11679 10655 11685
rect 10597 11645 10609 11679
rect 10643 11645 10655 11679
rect 10597 11639 10655 11645
rect 10781 11679 10839 11685
rect 10781 11645 10793 11679
rect 10827 11645 10839 11679
rect 10781 11639 10839 11645
rect 3234 11568 3240 11620
rect 3292 11608 3298 11620
rect 7006 11608 7012 11620
rect 3292 11580 7012 11608
rect 3292 11568 3298 11580
rect 7006 11568 7012 11580
rect 7064 11568 7070 11620
rect 7944 11608 7972 11636
rect 8573 11611 8631 11617
rect 8573 11608 8585 11611
rect 7944 11580 8585 11608
rect 8573 11577 8585 11580
rect 8619 11577 8631 11611
rect 8573 11571 8631 11577
rect 10321 11611 10379 11617
rect 10321 11577 10333 11611
rect 10367 11608 10379 11611
rect 10612 11608 10640 11639
rect 10367 11580 10640 11608
rect 10367 11577 10379 11580
rect 10321 11571 10379 11577
rect 10686 11568 10692 11620
rect 10744 11608 10750 11620
rect 10796 11608 10824 11639
rect 10870 11636 10876 11688
rect 10928 11636 10934 11688
rect 13078 11636 13084 11688
rect 13136 11676 13142 11688
rect 14654 11679 14712 11685
rect 14654 11676 14666 11679
rect 13136 11648 14666 11676
rect 13136 11636 13142 11648
rect 14654 11645 14666 11648
rect 14700 11645 14712 11679
rect 14654 11639 14712 11645
rect 15654 11636 15660 11688
rect 15712 11676 15718 11688
rect 16025 11679 16083 11685
rect 16025 11676 16037 11679
rect 15712 11648 16037 11676
rect 15712 11636 15718 11648
rect 16025 11645 16037 11648
rect 16071 11645 16083 11679
rect 16025 11639 16083 11645
rect 15010 11608 15016 11620
rect 10744 11580 15016 11608
rect 10744 11568 10750 11580
rect 15010 11568 15016 11580
rect 15068 11568 15074 11620
rect 16040 11608 16068 11639
rect 16114 11636 16120 11688
rect 16172 11676 16178 11688
rect 16485 11679 16543 11685
rect 16485 11676 16497 11679
rect 16172 11648 16497 11676
rect 16172 11636 16178 11648
rect 16485 11645 16497 11648
rect 16531 11645 16543 11679
rect 16485 11639 16543 11645
rect 16577 11679 16635 11685
rect 16577 11645 16589 11679
rect 16623 11645 16635 11679
rect 16577 11639 16635 11645
rect 16592 11608 16620 11639
rect 17310 11636 17316 11688
rect 17368 11636 17374 11688
rect 17512 11685 17540 11716
rect 17497 11679 17555 11685
rect 17497 11645 17509 11679
rect 17543 11645 17555 11679
rect 17497 11639 17555 11645
rect 19429 11679 19487 11685
rect 19429 11645 19441 11679
rect 19475 11645 19487 11679
rect 19429 11639 19487 11645
rect 19613 11679 19671 11685
rect 19613 11645 19625 11679
rect 19659 11676 19671 11679
rect 19889 11679 19947 11685
rect 19889 11676 19901 11679
rect 19659 11648 19901 11676
rect 19659 11645 19671 11648
rect 19613 11639 19671 11645
rect 19889 11645 19901 11648
rect 19935 11676 19947 11679
rect 20180 11676 20208 11775
rect 21560 11753 21588 11852
rect 21634 11840 21640 11892
rect 21692 11840 21698 11892
rect 21545 11747 21603 11753
rect 21545 11713 21557 11747
rect 21591 11713 21603 11747
rect 21545 11707 21603 11713
rect 19935 11648 20208 11676
rect 19935 11645 19947 11648
rect 19889 11639 19947 11645
rect 16040 11580 16620 11608
rect 19444 11608 19472 11639
rect 20714 11636 20720 11688
rect 20772 11676 20778 11688
rect 21278 11679 21336 11685
rect 21278 11676 21290 11679
rect 20772 11648 21290 11676
rect 20772 11636 20778 11648
rect 21278 11645 21290 11648
rect 21324 11645 21336 11679
rect 21560 11676 21588 11707
rect 22370 11676 22376 11688
rect 21560 11648 22376 11676
rect 21278 11639 21336 11645
rect 22370 11636 22376 11648
rect 22428 11676 22434 11688
rect 23017 11679 23075 11685
rect 23017 11676 23029 11679
rect 22428 11648 23029 11676
rect 22428 11636 22434 11648
rect 23017 11645 23029 11648
rect 23063 11645 23075 11679
rect 23017 11639 23075 11645
rect 19518 11608 19524 11620
rect 19444 11580 19524 11608
rect 19518 11568 19524 11580
rect 19576 11608 19582 11620
rect 19705 11611 19763 11617
rect 19705 11608 19717 11611
rect 19576 11580 19717 11608
rect 19576 11568 19582 11580
rect 19705 11577 19717 11580
rect 19751 11577 19763 11611
rect 19705 11571 19763 11577
rect 21818 11568 21824 11620
rect 21876 11608 21882 11620
rect 22750 11611 22808 11617
rect 22750 11608 22762 11611
rect 21876 11580 22762 11608
rect 21876 11568 21882 11580
rect 22750 11577 22762 11580
rect 22796 11577 22808 11611
rect 22750 11571 22808 11577
rect 4706 11500 4712 11552
rect 4764 11500 4770 11552
rect 5074 11500 5080 11552
rect 5132 11500 5138 11552
rect 8018 11500 8024 11552
rect 8076 11500 8082 11552
rect 8754 11500 8760 11552
rect 8812 11500 8818 11552
rect 9122 11500 9128 11552
rect 9180 11500 9186 11552
rect 10410 11500 10416 11552
rect 10468 11500 10474 11552
rect 13541 11543 13599 11549
rect 13541 11509 13553 11543
rect 13587 11540 13599 11543
rect 13630 11540 13636 11552
rect 13587 11512 13636 11540
rect 13587 11509 13599 11512
rect 13541 11503 13599 11509
rect 13630 11500 13636 11512
rect 13688 11500 13694 11552
rect 552 11450 23368 11472
rect 552 11398 4322 11450
rect 4374 11398 4386 11450
rect 4438 11398 4450 11450
rect 4502 11398 4514 11450
rect 4566 11398 4578 11450
rect 4630 11398 23368 11450
rect 552 11376 23368 11398
rect 4617 11339 4675 11345
rect 4617 11305 4629 11339
rect 4663 11336 4675 11339
rect 5074 11336 5080 11348
rect 4663 11308 5080 11336
rect 4663 11305 4675 11308
rect 4617 11299 4675 11305
rect 5074 11296 5080 11308
rect 5132 11296 5138 11348
rect 6178 11296 6184 11348
rect 6236 11336 6242 11348
rect 6273 11339 6331 11345
rect 6273 11336 6285 11339
rect 6236 11308 6285 11336
rect 6236 11296 6242 11308
rect 6273 11305 6285 11308
rect 6319 11305 6331 11339
rect 6273 11299 6331 11305
rect 10781 11339 10839 11345
rect 10781 11305 10793 11339
rect 10827 11336 10839 11339
rect 10870 11336 10876 11348
rect 10827 11308 10876 11336
rect 10827 11305 10839 11308
rect 10781 11299 10839 11305
rect 10870 11296 10876 11308
rect 10928 11296 10934 11348
rect 11333 11339 11391 11345
rect 11333 11305 11345 11339
rect 11379 11336 11391 11339
rect 12250 11336 12256 11348
rect 11379 11308 12256 11336
rect 11379 11305 11391 11308
rect 11333 11299 11391 11305
rect 3504 11271 3562 11277
rect 3504 11237 3516 11271
rect 3550 11268 3562 11271
rect 4706 11268 4712 11280
rect 3550 11240 4712 11268
rect 3550 11237 3562 11240
rect 3504 11231 3562 11237
rect 4706 11228 4712 11240
rect 4764 11228 4770 11280
rect 7006 11228 7012 11280
rect 7064 11268 7070 11280
rect 11348 11268 11376 11299
rect 12250 11296 12256 11308
rect 12308 11296 12314 11348
rect 13538 11296 13544 11348
rect 13596 11296 13602 11348
rect 18046 11296 18052 11348
rect 18104 11336 18110 11348
rect 18433 11339 18491 11345
rect 18433 11336 18445 11339
rect 18104 11308 18445 11336
rect 18104 11296 18110 11308
rect 18433 11305 18445 11308
rect 18479 11305 18491 11339
rect 18433 11299 18491 11305
rect 21818 11296 21824 11348
rect 21876 11296 21882 11348
rect 7064 11240 11376 11268
rect 7064 11228 7070 11240
rect 6181 11203 6239 11209
rect 6181 11169 6193 11203
rect 6227 11200 6239 11203
rect 6730 11200 6736 11212
rect 6227 11172 6736 11200
rect 6227 11169 6239 11172
rect 6181 11163 6239 11169
rect 6730 11160 6736 11172
rect 6788 11160 6794 11212
rect 8018 11160 8024 11212
rect 8076 11160 8082 11212
rect 8205 11203 8263 11209
rect 8205 11169 8217 11203
rect 8251 11200 8263 11203
rect 8754 11200 8760 11212
rect 8251 11172 8760 11200
rect 8251 11169 8263 11172
rect 8205 11163 8263 11169
rect 8754 11160 8760 11172
rect 8812 11160 8818 11212
rect 10502 11160 10508 11212
rect 10560 11160 10566 11212
rect 10612 11209 10640 11240
rect 18138 11228 18144 11280
rect 18196 11268 18202 11280
rect 18233 11271 18291 11277
rect 18233 11268 18245 11271
rect 18196 11240 18245 11268
rect 18196 11228 18202 11240
rect 18233 11237 18245 11240
rect 18279 11237 18291 11271
rect 18233 11231 18291 11237
rect 19334 11228 19340 11280
rect 19392 11268 19398 11280
rect 19889 11271 19947 11277
rect 19889 11268 19901 11271
rect 19392 11240 19901 11268
rect 19392 11228 19398 11240
rect 19889 11237 19901 11240
rect 19935 11268 19947 11271
rect 20622 11268 20628 11280
rect 19935 11240 20628 11268
rect 19935 11237 19947 11240
rect 19889 11231 19947 11237
rect 20622 11228 20628 11240
rect 20680 11228 20686 11280
rect 21542 11228 21548 11280
rect 21600 11268 21606 11280
rect 21637 11271 21695 11277
rect 21637 11268 21649 11271
rect 21600 11240 21649 11268
rect 21600 11228 21606 11240
rect 21637 11237 21649 11240
rect 21683 11237 21695 11271
rect 21637 11231 21695 11237
rect 22002 11228 22008 11280
rect 22060 11228 22066 11280
rect 10597 11203 10655 11209
rect 10597 11169 10609 11203
rect 10643 11169 10655 11203
rect 10597 11163 10655 11169
rect 11238 11160 11244 11212
rect 11296 11160 11302 11212
rect 11698 11160 11704 11212
rect 11756 11160 11762 11212
rect 11793 11203 11851 11209
rect 11793 11169 11805 11203
rect 11839 11200 11851 11203
rect 12434 11200 12440 11212
rect 11839 11172 12440 11200
rect 11839 11169 11851 11172
rect 11793 11163 11851 11169
rect 12434 11160 12440 11172
rect 12492 11160 12498 11212
rect 13725 11203 13783 11209
rect 13725 11169 13737 11203
rect 13771 11200 13783 11203
rect 15470 11200 15476 11212
rect 13771 11172 15476 11200
rect 13771 11169 13783 11172
rect 13725 11163 13783 11169
rect 15470 11160 15476 11172
rect 15528 11160 15534 11212
rect 15565 11203 15623 11209
rect 15565 11169 15577 11203
rect 15611 11200 15623 11203
rect 16114 11200 16120 11212
rect 15611 11172 16120 11200
rect 15611 11169 15623 11172
rect 15565 11163 15623 11169
rect 16114 11160 16120 11172
rect 16172 11160 16178 11212
rect 19150 11160 19156 11212
rect 19208 11200 19214 11212
rect 19429 11203 19487 11209
rect 19429 11200 19441 11203
rect 19208 11172 19441 11200
rect 19208 11160 19214 11172
rect 19429 11169 19441 11172
rect 19475 11169 19487 11203
rect 19429 11163 19487 11169
rect 20073 11203 20131 11209
rect 20073 11169 20085 11203
rect 20119 11200 20131 11203
rect 20809 11203 20867 11209
rect 20809 11200 20821 11203
rect 20119 11172 20821 11200
rect 20119 11169 20131 11172
rect 20073 11163 20131 11169
rect 20809 11169 20821 11172
rect 20855 11169 20867 11203
rect 20809 11163 20867 11169
rect 3234 11092 3240 11144
rect 3292 11092 3298 11144
rect 5258 11092 5264 11144
rect 5316 11132 5322 11144
rect 6365 11135 6423 11141
rect 6365 11132 6377 11135
rect 5316 11104 6377 11132
rect 5316 11092 5322 11104
rect 6365 11101 6377 11104
rect 6411 11132 6423 11135
rect 10686 11132 10692 11144
rect 6411 11104 10692 11132
rect 6411 11101 6423 11104
rect 6365 11095 6423 11101
rect 10686 11092 10692 11104
rect 10744 11092 10750 11144
rect 12894 11092 12900 11144
rect 12952 11132 12958 11144
rect 13630 11132 13636 11144
rect 12952 11104 13636 11132
rect 12952 11092 12958 11104
rect 13630 11092 13636 11104
rect 13688 11132 13694 11144
rect 13909 11135 13967 11141
rect 13909 11132 13921 11135
rect 13688 11104 13921 11132
rect 13688 11092 13694 11104
rect 13909 11101 13921 11104
rect 13955 11101 13967 11135
rect 13909 11095 13967 11101
rect 15654 11092 15660 11144
rect 15712 11092 15718 11144
rect 19245 11135 19303 11141
rect 19245 11101 19257 11135
rect 19291 11132 19303 11135
rect 19334 11132 19340 11144
rect 19291 11104 19340 11132
rect 19291 11101 19303 11104
rect 19245 11095 19303 11101
rect 19334 11092 19340 11104
rect 19392 11092 19398 11144
rect 19444 11132 19472 11163
rect 20088 11132 20116 11163
rect 19444 11104 20116 11132
rect 20533 11135 20591 11141
rect 20533 11101 20545 11135
rect 20579 11101 20591 11135
rect 20533 11095 20591 11101
rect 20548 11064 20576 11095
rect 20622 11092 20628 11144
rect 20680 11092 20686 11144
rect 20714 11092 20720 11144
rect 20772 11092 20778 11144
rect 20806 11064 20812 11076
rect 20548 11036 20812 11064
rect 20806 11024 20812 11036
rect 20864 11024 20870 11076
rect 20898 11024 20904 11076
rect 20956 11064 20962 11076
rect 21269 11067 21327 11073
rect 21269 11064 21281 11067
rect 20956 11036 21281 11064
rect 20956 11024 20962 11036
rect 21269 11033 21281 11036
rect 21315 11033 21327 11067
rect 21269 11027 21327 11033
rect 22094 11024 22100 11076
rect 22152 11064 22158 11076
rect 22189 11067 22247 11073
rect 22189 11064 22201 11067
rect 22152 11036 22201 11064
rect 22152 11024 22158 11036
rect 22189 11033 22201 11036
rect 22235 11033 22247 11067
rect 22189 11027 22247 11033
rect 5626 10956 5632 11008
rect 5684 10996 5690 11008
rect 5813 10999 5871 11005
rect 5813 10996 5825 10999
rect 5684 10968 5825 10996
rect 5684 10956 5690 10968
rect 5813 10965 5825 10968
rect 5859 10965 5871 10999
rect 5813 10959 5871 10965
rect 8110 10956 8116 11008
rect 8168 10956 8174 11008
rect 11606 10956 11612 11008
rect 11664 10956 11670 11008
rect 15930 10956 15936 11008
rect 15988 10956 15994 11008
rect 18414 10956 18420 11008
rect 18472 10956 18478 11008
rect 18601 10999 18659 11005
rect 18601 10965 18613 10999
rect 18647 10996 18659 10999
rect 19150 10996 19156 11008
rect 18647 10968 19156 10996
rect 18647 10965 18659 10968
rect 18601 10959 18659 10965
rect 19150 10956 19156 10968
rect 19208 10956 19214 11008
rect 19518 10956 19524 11008
rect 19576 10996 19582 11008
rect 19613 10999 19671 11005
rect 19613 10996 19625 10999
rect 19576 10968 19625 10996
rect 19576 10956 19582 10968
rect 19613 10965 19625 10968
rect 19659 10965 19671 10999
rect 19613 10959 19671 10965
rect 19705 10999 19763 11005
rect 19705 10965 19717 10999
rect 19751 10996 19763 10999
rect 19886 10996 19892 11008
rect 19751 10968 19892 10996
rect 19751 10965 19763 10968
rect 19705 10959 19763 10965
rect 19886 10956 19892 10968
rect 19944 10956 19950 11008
rect 20993 10999 21051 11005
rect 20993 10965 21005 10999
rect 21039 10996 21051 10999
rect 21637 10999 21695 11005
rect 21637 10996 21649 10999
rect 21039 10968 21649 10996
rect 21039 10965 21051 10968
rect 20993 10959 21051 10965
rect 21637 10965 21649 10968
rect 21683 10965 21695 10999
rect 21637 10959 21695 10965
rect 552 10906 23368 10928
rect 552 10854 3662 10906
rect 3714 10854 3726 10906
rect 3778 10854 3790 10906
rect 3842 10854 3854 10906
rect 3906 10854 3918 10906
rect 3970 10854 23368 10906
rect 552 10832 23368 10854
rect 6730 10752 6736 10804
rect 6788 10752 6794 10804
rect 8110 10752 8116 10804
rect 8168 10792 8174 10804
rect 8481 10795 8539 10801
rect 8481 10792 8493 10795
rect 8168 10764 8493 10792
rect 8168 10752 8174 10764
rect 8481 10761 8493 10764
rect 8527 10761 8539 10795
rect 8481 10755 8539 10761
rect 10502 10752 10508 10804
rect 10560 10792 10566 10804
rect 10962 10792 10968 10804
rect 10560 10764 10968 10792
rect 10560 10752 10566 10764
rect 10962 10752 10968 10764
rect 11020 10752 11026 10804
rect 11238 10752 11244 10804
rect 11296 10792 11302 10804
rect 12437 10795 12495 10801
rect 12437 10792 12449 10795
rect 11296 10764 12449 10792
rect 11296 10752 11302 10764
rect 12437 10761 12449 10764
rect 12483 10761 12495 10795
rect 12437 10755 12495 10761
rect 18506 10752 18512 10804
rect 18564 10792 18570 10804
rect 18877 10795 18935 10801
rect 18877 10792 18889 10795
rect 18564 10764 18889 10792
rect 18564 10752 18570 10764
rect 18877 10761 18889 10764
rect 18923 10761 18935 10795
rect 18877 10755 18935 10761
rect 19334 10752 19340 10804
rect 19392 10752 19398 10804
rect 20806 10752 20812 10804
rect 20864 10792 20870 10804
rect 20993 10795 21051 10801
rect 20993 10792 21005 10795
rect 20864 10764 21005 10792
rect 20864 10752 20870 10764
rect 20993 10761 21005 10764
rect 21039 10792 21051 10795
rect 21634 10792 21640 10804
rect 21039 10764 21640 10792
rect 21039 10761 21051 10764
rect 20993 10755 21051 10761
rect 21634 10752 21640 10764
rect 21692 10752 21698 10804
rect 7929 10659 7987 10665
rect 7929 10625 7941 10659
rect 7975 10656 7987 10659
rect 8128 10656 8156 10752
rect 19150 10684 19156 10736
rect 19208 10724 19214 10736
rect 19245 10727 19303 10733
rect 19245 10724 19257 10727
rect 19208 10696 19257 10724
rect 19208 10684 19214 10696
rect 19245 10693 19257 10696
rect 19291 10693 19303 10727
rect 19245 10687 19303 10693
rect 20898 10684 20904 10736
rect 20956 10724 20962 10736
rect 21177 10727 21235 10733
rect 21177 10724 21189 10727
rect 20956 10696 21189 10724
rect 20956 10684 20962 10696
rect 21177 10693 21189 10696
rect 21223 10693 21235 10727
rect 21177 10687 21235 10693
rect 7975 10628 8156 10656
rect 8849 10659 8907 10665
rect 7975 10625 7987 10628
rect 7929 10619 7987 10625
rect 8849 10625 8861 10659
rect 8895 10656 8907 10659
rect 9033 10659 9091 10665
rect 9033 10656 9045 10659
rect 8895 10628 9045 10656
rect 8895 10625 8907 10628
rect 8849 10619 8907 10625
rect 9033 10625 9045 10628
rect 9079 10625 9091 10659
rect 9033 10619 9091 10625
rect 14090 10616 14096 10668
rect 14148 10616 14154 10668
rect 14274 10616 14280 10668
rect 14332 10656 14338 10668
rect 14550 10656 14556 10668
rect 14332 10628 14556 10656
rect 14332 10616 14338 10628
rect 14550 10616 14556 10628
rect 14608 10616 14614 10668
rect 5350 10548 5356 10600
rect 5408 10548 5414 10600
rect 5626 10597 5632 10600
rect 5620 10588 5632 10597
rect 5587 10560 5632 10588
rect 5620 10551 5632 10560
rect 5626 10548 5632 10551
rect 5684 10548 5690 10600
rect 7006 10548 7012 10600
rect 7064 10588 7070 10600
rect 7193 10591 7251 10597
rect 7193 10588 7205 10591
rect 7064 10560 7205 10588
rect 7064 10548 7070 10560
rect 7193 10557 7205 10560
rect 7239 10557 7251 10591
rect 7193 10551 7251 10557
rect 7558 10548 7564 10600
rect 7616 10548 7622 10600
rect 7834 10548 7840 10600
rect 7892 10548 7898 10600
rect 8389 10591 8447 10597
rect 8389 10557 8401 10591
rect 8435 10557 8447 10591
rect 8389 10551 8447 10557
rect 8665 10591 8723 10597
rect 8665 10557 8677 10591
rect 8711 10588 8723 10591
rect 8754 10588 8760 10600
rect 8711 10560 8760 10588
rect 8711 10557 8723 10560
rect 8665 10551 8723 10557
rect 7282 10480 7288 10532
rect 7340 10480 7346 10532
rect 7377 10523 7435 10529
rect 7377 10489 7389 10523
rect 7423 10520 7435 10523
rect 8110 10520 8116 10532
rect 7423 10492 8116 10520
rect 7423 10489 7435 10492
rect 7377 10483 7435 10489
rect 8110 10480 8116 10492
rect 8168 10520 8174 10532
rect 8404 10520 8432 10551
rect 8754 10548 8760 10560
rect 8812 10548 8818 10600
rect 9122 10548 9128 10600
rect 9180 10548 9186 10600
rect 9585 10591 9643 10597
rect 9585 10557 9597 10591
rect 9631 10557 9643 10591
rect 9585 10551 9643 10557
rect 9852 10591 9910 10597
rect 9852 10557 9864 10591
rect 9898 10588 9910 10591
rect 10410 10588 10416 10600
rect 9898 10560 10416 10588
rect 9898 10557 9910 10560
rect 9852 10551 9910 10557
rect 8168 10492 8432 10520
rect 8168 10480 8174 10492
rect 9398 10480 9404 10532
rect 9456 10520 9462 10532
rect 9600 10520 9628 10551
rect 10410 10548 10416 10560
rect 10468 10548 10474 10600
rect 11057 10591 11115 10597
rect 11057 10557 11069 10591
rect 11103 10557 11115 10591
rect 11057 10551 11115 10557
rect 11324 10591 11382 10597
rect 11324 10557 11336 10591
rect 11370 10588 11382 10591
rect 11606 10588 11612 10600
rect 11370 10560 11612 10588
rect 11370 10557 11382 10560
rect 11324 10551 11382 10557
rect 11072 10520 11100 10551
rect 11606 10548 11612 10560
rect 11664 10548 11670 10600
rect 18509 10591 18567 10597
rect 18509 10557 18521 10591
rect 18555 10588 18567 10591
rect 19242 10588 19248 10600
rect 18555 10560 19248 10588
rect 18555 10557 18567 10560
rect 18509 10551 18567 10557
rect 19242 10548 19248 10560
rect 19300 10588 19306 10600
rect 20717 10591 20775 10597
rect 20717 10588 20729 10591
rect 19300 10560 20729 10588
rect 19300 10548 19306 10560
rect 20717 10557 20729 10560
rect 20763 10588 20775 10591
rect 21174 10588 21180 10600
rect 20763 10560 21180 10588
rect 20763 10557 20775 10560
rect 20717 10551 20775 10557
rect 21174 10548 21180 10560
rect 21232 10548 21238 10600
rect 9456 10492 11100 10520
rect 18264 10523 18322 10529
rect 9456 10480 9462 10492
rect 18264 10489 18276 10523
rect 18310 10520 18322 10523
rect 18310 10492 18736 10520
rect 18310 10489 18322 10492
rect 18264 10483 18322 10489
rect 7006 10412 7012 10464
rect 7064 10412 7070 10464
rect 8205 10455 8263 10461
rect 8205 10421 8217 10455
rect 8251 10452 8263 10455
rect 8846 10452 8852 10464
rect 8251 10424 8852 10452
rect 8251 10421 8263 10424
rect 8205 10415 8263 10421
rect 8846 10412 8852 10424
rect 8904 10412 8910 10464
rect 9493 10455 9551 10461
rect 9493 10421 9505 10455
rect 9539 10452 9551 10455
rect 10502 10452 10508 10464
rect 9539 10424 10508 10452
rect 9539 10421 9551 10424
rect 9493 10415 9551 10421
rect 10502 10412 10508 10424
rect 10560 10412 10566 10464
rect 13633 10455 13691 10461
rect 13633 10421 13645 10455
rect 13679 10452 13691 10455
rect 13814 10452 13820 10464
rect 13679 10424 13820 10452
rect 13679 10421 13691 10424
rect 13633 10415 13691 10421
rect 13814 10412 13820 10424
rect 13872 10412 13878 10464
rect 13906 10412 13912 10464
rect 13964 10452 13970 10464
rect 14001 10455 14059 10461
rect 14001 10452 14013 10455
rect 13964 10424 14013 10452
rect 13964 10412 13970 10424
rect 14001 10421 14013 10424
rect 14047 10421 14059 10455
rect 14001 10415 14059 10421
rect 17129 10455 17187 10461
rect 17129 10421 17141 10455
rect 17175 10452 17187 10455
rect 18414 10452 18420 10464
rect 17175 10424 18420 10452
rect 17175 10421 17187 10424
rect 17129 10415 17187 10421
rect 18414 10412 18420 10424
rect 18472 10412 18478 10464
rect 18708 10461 18736 10492
rect 20070 10480 20076 10532
rect 20128 10520 20134 10532
rect 20450 10523 20508 10529
rect 20450 10520 20462 10523
rect 20128 10492 20462 10520
rect 20128 10480 20134 10492
rect 20450 10489 20462 10492
rect 20496 10489 20508 10523
rect 20450 10483 20508 10489
rect 20806 10480 20812 10532
rect 20864 10480 20870 10532
rect 18693 10455 18751 10461
rect 18693 10421 18705 10455
rect 18739 10421 18751 10455
rect 18693 10415 18751 10421
rect 18874 10412 18880 10464
rect 18932 10412 18938 10464
rect 19518 10412 19524 10464
rect 19576 10452 19582 10464
rect 21009 10455 21067 10461
rect 21009 10452 21021 10455
rect 19576 10424 21021 10452
rect 19576 10412 19582 10424
rect 21009 10421 21021 10424
rect 21055 10421 21067 10455
rect 21009 10415 21067 10421
rect 552 10362 23368 10384
rect 552 10310 4322 10362
rect 4374 10310 4386 10362
rect 4438 10310 4450 10362
rect 4502 10310 4514 10362
rect 4566 10310 4578 10362
rect 4630 10310 23368 10362
rect 552 10288 23368 10310
rect 4709 10251 4767 10257
rect 4709 10217 4721 10251
rect 4755 10248 4767 10251
rect 5442 10248 5448 10260
rect 4755 10220 5448 10248
rect 4755 10217 4767 10220
rect 4709 10211 4767 10217
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 7282 10208 7288 10260
rect 7340 10248 7346 10260
rect 7742 10248 7748 10260
rect 7340 10220 7748 10248
rect 7340 10208 7346 10220
rect 7742 10208 7748 10220
rect 7800 10248 7806 10260
rect 7929 10251 7987 10257
rect 7929 10248 7941 10251
rect 7800 10220 7941 10248
rect 7800 10208 7806 10220
rect 7929 10217 7941 10220
rect 7975 10217 7987 10251
rect 7929 10211 7987 10217
rect 8110 10208 8116 10260
rect 8168 10208 8174 10260
rect 16669 10251 16727 10257
rect 16669 10217 16681 10251
rect 16715 10217 16727 10251
rect 16669 10211 16727 10217
rect 17221 10251 17279 10257
rect 17221 10217 17233 10251
rect 17267 10248 17279 10251
rect 17954 10248 17960 10260
rect 17267 10220 17960 10248
rect 17267 10217 17279 10220
rect 17221 10211 17279 10217
rect 6816 10183 6874 10189
rect 4264 10152 4844 10180
rect 3326 10072 3332 10124
rect 3384 10112 3390 10124
rect 3384 10084 3832 10112
rect 3384 10072 3390 10084
rect 3421 10047 3479 10053
rect 3421 10013 3433 10047
rect 3467 10044 3479 10047
rect 3510 10044 3516 10056
rect 3467 10016 3516 10044
rect 3467 10013 3479 10016
rect 3421 10007 3479 10013
rect 3510 10004 3516 10016
rect 3568 10004 3574 10056
rect 3804 10044 3832 10084
rect 4264 10044 4292 10152
rect 4816 10121 4844 10152
rect 6816 10149 6828 10183
rect 6862 10180 6874 10183
rect 7006 10180 7012 10192
rect 6862 10152 7012 10180
rect 6862 10149 6874 10152
rect 6816 10143 6874 10149
rect 7006 10140 7012 10152
rect 7064 10140 7070 10192
rect 13848 10183 13906 10189
rect 13848 10149 13860 10183
rect 13894 10180 13906 10183
rect 14185 10183 14243 10189
rect 14185 10180 14197 10183
rect 13894 10152 14197 10180
rect 13894 10149 13906 10152
rect 13848 10143 13906 10149
rect 14185 10149 14197 10152
rect 14231 10149 14243 10183
rect 14185 10143 14243 10149
rect 15565 10183 15623 10189
rect 15565 10149 15577 10183
rect 15611 10149 15623 10183
rect 15565 10143 15623 10149
rect 4341 10115 4399 10121
rect 4341 10081 4353 10115
rect 4387 10112 4399 10115
rect 4801 10115 4859 10121
rect 4387 10084 4752 10112
rect 4387 10081 4399 10084
rect 4341 10075 4399 10081
rect 4724 10056 4752 10084
rect 4801 10081 4813 10115
rect 4847 10112 4859 10115
rect 4890 10112 4896 10124
rect 4847 10084 4896 10112
rect 4847 10081 4859 10084
rect 4801 10075 4859 10081
rect 4890 10072 4896 10084
rect 4948 10072 4954 10124
rect 5350 10072 5356 10124
rect 5408 10112 5414 10124
rect 6549 10115 6607 10121
rect 6549 10112 6561 10115
rect 5408 10084 6561 10112
rect 5408 10072 5414 10084
rect 6549 10081 6561 10084
rect 6595 10112 6607 10115
rect 6595 10084 7788 10112
rect 6595 10081 6607 10084
rect 6549 10075 6607 10081
rect 4433 10047 4491 10053
rect 4433 10044 4445 10047
rect 3804 10016 4445 10044
rect 4433 10013 4445 10016
rect 4479 10013 4491 10047
rect 4433 10007 4491 10013
rect 4706 10004 4712 10056
rect 4764 10044 4770 10056
rect 5074 10044 5080 10056
rect 4764 10016 5080 10044
rect 4764 10004 4770 10016
rect 5074 10004 5080 10016
rect 5132 10004 5138 10056
rect 7760 10044 7788 10084
rect 7834 10072 7840 10124
rect 7892 10112 7898 10124
rect 8021 10115 8079 10121
rect 8021 10112 8033 10115
rect 7892 10084 8033 10112
rect 7892 10072 7898 10084
rect 8021 10081 8033 10084
rect 8067 10081 8079 10115
rect 8021 10075 8079 10081
rect 13998 10072 14004 10124
rect 14056 10112 14062 10124
rect 14093 10115 14151 10121
rect 14093 10112 14105 10115
rect 14056 10084 14105 10112
rect 14056 10072 14062 10084
rect 14093 10081 14105 10084
rect 14139 10081 14151 10115
rect 14093 10075 14151 10081
rect 14366 10072 14372 10124
rect 14424 10072 14430 10124
rect 14550 10072 14556 10124
rect 14608 10072 14614 10124
rect 9398 10044 9404 10056
rect 7760 10016 9404 10044
rect 9398 10004 9404 10016
rect 9456 10004 9462 10056
rect 14645 10047 14703 10053
rect 14645 10013 14657 10047
rect 14691 10013 14703 10047
rect 15580 10044 15608 10143
rect 15746 10140 15752 10192
rect 15804 10189 15810 10192
rect 15804 10183 15823 10189
rect 15811 10149 15823 10183
rect 16684 10180 16712 10211
rect 17954 10208 17960 10220
rect 18012 10208 18018 10260
rect 18138 10208 18144 10260
rect 18196 10208 18202 10260
rect 18506 10208 18512 10260
rect 18564 10208 18570 10260
rect 20070 10208 20076 10260
rect 20128 10208 20134 10260
rect 20898 10208 20904 10260
rect 20956 10248 20962 10260
rect 22071 10251 22129 10257
rect 22071 10248 22083 10251
rect 20956 10220 22083 10248
rect 20956 10208 20962 10220
rect 22071 10217 22083 10220
rect 22117 10217 22129 10251
rect 22071 10211 22129 10217
rect 16684 10152 17080 10180
rect 15804 10143 15823 10149
rect 15804 10140 15810 10143
rect 16301 10115 16359 10121
rect 16301 10081 16313 10115
rect 16347 10112 16359 10115
rect 16574 10112 16580 10124
rect 16347 10084 16580 10112
rect 16347 10081 16359 10084
rect 16301 10075 16359 10081
rect 16574 10072 16580 10084
rect 16632 10072 16638 10124
rect 16758 10072 16764 10124
rect 16816 10072 16822 10124
rect 17052 10121 17080 10152
rect 18874 10140 18880 10192
rect 18932 10180 18938 10192
rect 19889 10183 19947 10189
rect 19889 10180 19901 10183
rect 18932 10152 19901 10180
rect 18932 10140 18938 10152
rect 19889 10149 19901 10152
rect 19935 10180 19947 10183
rect 20990 10180 20996 10192
rect 19935 10152 20996 10180
rect 19935 10149 19947 10152
rect 19889 10143 19947 10149
rect 20990 10140 20996 10152
rect 21048 10140 21054 10192
rect 21453 10183 21511 10189
rect 21453 10149 21465 10183
rect 21499 10180 21511 10183
rect 21542 10180 21548 10192
rect 21499 10152 21548 10180
rect 21499 10149 21511 10152
rect 21453 10143 21511 10149
rect 17037 10115 17095 10121
rect 17037 10081 17049 10115
rect 17083 10081 17095 10115
rect 17037 10075 17095 10081
rect 18046 10072 18052 10124
rect 18104 10072 18110 10124
rect 18325 10115 18383 10121
rect 18325 10081 18337 10115
rect 18371 10112 18383 10115
rect 18414 10112 18420 10124
rect 18371 10084 18420 10112
rect 18371 10081 18383 10084
rect 18325 10075 18383 10081
rect 18414 10072 18420 10084
rect 18472 10072 18478 10124
rect 19518 10072 19524 10124
rect 19576 10072 19582 10124
rect 20714 10072 20720 10124
rect 20772 10112 20778 10124
rect 21468 10112 21496 10143
rect 21542 10140 21548 10152
rect 21600 10140 21606 10192
rect 22186 10140 22192 10192
rect 22244 10180 22250 10192
rect 22281 10183 22339 10189
rect 22281 10180 22293 10183
rect 22244 10152 22293 10180
rect 22244 10140 22250 10152
rect 22281 10149 22293 10152
rect 22327 10180 22339 10183
rect 22462 10180 22468 10192
rect 22327 10152 22468 10180
rect 22327 10149 22339 10152
rect 22281 10143 22339 10149
rect 22462 10140 22468 10152
rect 22520 10140 22526 10192
rect 22554 10140 22560 10192
rect 22612 10140 22618 10192
rect 22373 10115 22431 10121
rect 22373 10112 22385 10115
rect 20772 10084 21496 10112
rect 21836 10084 22385 10112
rect 20772 10072 20778 10084
rect 15838 10044 15844 10056
rect 15580 10016 15844 10044
rect 14645 10007 14703 10013
rect 3528 9976 3556 10004
rect 3528 9948 4384 9976
rect 3697 9911 3755 9917
rect 3697 9877 3709 9911
rect 3743 9908 3755 9911
rect 4062 9908 4068 9920
rect 3743 9880 4068 9908
rect 3743 9877 3755 9880
rect 3697 9871 3755 9877
rect 4062 9868 4068 9880
rect 4120 9868 4126 9920
rect 4356 9917 4384 9948
rect 4798 9936 4804 9988
rect 4856 9976 4862 9988
rect 4985 9979 5043 9985
rect 4985 9976 4997 9979
rect 4856 9948 4997 9976
rect 4856 9936 4862 9948
rect 4985 9945 4997 9948
rect 5031 9945 5043 9979
rect 4985 9939 5043 9945
rect 4341 9911 4399 9917
rect 4341 9877 4353 9911
rect 4387 9908 4399 9911
rect 4614 9908 4620 9920
rect 4387 9880 4620 9908
rect 4387 9877 4399 9880
rect 4341 9871 4399 9877
rect 4614 9868 4620 9880
rect 4672 9908 4678 9920
rect 4893 9911 4951 9917
rect 4893 9908 4905 9911
rect 4672 9880 4905 9908
rect 4672 9868 4678 9880
rect 4893 9877 4905 9880
rect 4939 9877 4951 9911
rect 4893 9871 4951 9877
rect 12710 9868 12716 9920
rect 12768 9908 12774 9920
rect 14182 9908 14188 9920
rect 12768 9880 14188 9908
rect 12768 9868 12774 9880
rect 14182 9868 14188 9880
rect 14240 9908 14246 9920
rect 14660 9908 14688 10007
rect 15838 10004 15844 10016
rect 15896 10004 15902 10056
rect 15930 10004 15936 10056
rect 15988 10044 15994 10056
rect 16209 10047 16267 10053
rect 16209 10044 16221 10047
rect 15988 10016 16221 10044
rect 15988 10004 15994 10016
rect 16209 10013 16221 10016
rect 16255 10013 16267 10047
rect 16209 10007 16267 10013
rect 16850 10004 16856 10056
rect 16908 10004 16914 10056
rect 15948 9948 16804 9976
rect 14240 9880 14688 9908
rect 14240 9868 14246 9880
rect 15654 9868 15660 9920
rect 15712 9908 15718 9920
rect 15948 9917 15976 9948
rect 16776 9917 16804 9948
rect 20806 9936 20812 9988
rect 20864 9976 20870 9988
rect 21836 9985 21864 10084
rect 22373 10081 22385 10084
rect 22419 10081 22431 10115
rect 22373 10075 22431 10081
rect 21821 9979 21879 9985
rect 21821 9976 21833 9979
rect 20864 9948 21833 9976
rect 20864 9936 20870 9948
rect 21821 9945 21833 9948
rect 21867 9945 21879 9979
rect 21821 9939 21879 9945
rect 22002 9936 22008 9988
rect 22060 9976 22066 9988
rect 22741 9979 22799 9985
rect 22741 9976 22753 9979
rect 22060 9948 22753 9976
rect 22060 9936 22066 9948
rect 22741 9945 22753 9948
rect 22787 9945 22799 9979
rect 22741 9939 22799 9945
rect 15749 9911 15807 9917
rect 15749 9908 15761 9911
rect 15712 9880 15761 9908
rect 15712 9868 15718 9880
rect 15749 9877 15761 9880
rect 15795 9877 15807 9911
rect 15749 9871 15807 9877
rect 15933 9911 15991 9917
rect 15933 9877 15945 9911
rect 15979 9877 15991 9911
rect 15933 9871 15991 9877
rect 16761 9911 16819 9917
rect 16761 9877 16773 9911
rect 16807 9877 16819 9911
rect 16761 9871 16819 9877
rect 19886 9868 19892 9920
rect 19944 9868 19950 9920
rect 21266 9868 21272 9920
rect 21324 9868 21330 9920
rect 21358 9868 21364 9920
rect 21416 9908 21422 9920
rect 21453 9911 21511 9917
rect 21453 9908 21465 9911
rect 21416 9880 21465 9908
rect 21416 9868 21422 9880
rect 21453 9877 21465 9880
rect 21499 9877 21511 9911
rect 21453 9871 21511 9877
rect 21910 9868 21916 9920
rect 21968 9868 21974 9920
rect 22097 9911 22155 9917
rect 22097 9877 22109 9911
rect 22143 9908 22155 9911
rect 22554 9908 22560 9920
rect 22143 9880 22560 9908
rect 22143 9877 22155 9880
rect 22097 9871 22155 9877
rect 22554 9868 22560 9880
rect 22612 9868 22618 9920
rect 552 9818 23368 9840
rect 552 9766 3662 9818
rect 3714 9766 3726 9818
rect 3778 9766 3790 9818
rect 3842 9766 3854 9818
rect 3906 9766 3918 9818
rect 3970 9766 23368 9818
rect 552 9744 23368 9766
rect 4614 9664 4620 9716
rect 4672 9664 4678 9716
rect 5000 9676 5396 9704
rect 5000 9648 5028 9676
rect 4982 9636 4988 9648
rect 4632 9608 4988 9636
rect 4632 9509 4660 9608
rect 4982 9596 4988 9608
rect 5040 9596 5046 9648
rect 5074 9596 5080 9648
rect 5132 9636 5138 9648
rect 5261 9639 5319 9645
rect 5261 9636 5273 9639
rect 5132 9608 5273 9636
rect 5132 9596 5138 9608
rect 5261 9605 5273 9608
rect 5307 9605 5319 9639
rect 5368 9636 5396 9676
rect 12710 9664 12716 9716
rect 12768 9704 12774 9716
rect 13035 9707 13093 9713
rect 13035 9704 13047 9707
rect 12768 9676 13047 9704
rect 12768 9664 12774 9676
rect 13035 9673 13047 9676
rect 13081 9673 13093 9707
rect 13906 9704 13912 9716
rect 13035 9667 13093 9673
rect 13556 9676 13912 9704
rect 5368 9608 5764 9636
rect 5261 9599 5319 9605
rect 4706 9528 4712 9580
rect 4764 9528 4770 9580
rect 4798 9528 4804 9580
rect 4856 9568 4862 9580
rect 4856 9540 5580 9568
rect 4856 9528 4862 9540
rect 4617 9503 4675 9509
rect 4617 9469 4629 9503
rect 4663 9469 4675 9503
rect 4617 9463 4675 9469
rect 4890 9460 4896 9512
rect 4948 9460 4954 9512
rect 5442 9460 5448 9512
rect 5500 9460 5506 9512
rect 5552 9509 5580 9540
rect 5537 9503 5595 9509
rect 5537 9469 5549 9503
rect 5583 9469 5595 9503
rect 5537 9463 5595 9469
rect 5629 9503 5687 9509
rect 5629 9469 5641 9503
rect 5675 9469 5687 9503
rect 5736 9500 5764 9608
rect 9048 9608 10732 9636
rect 8846 9528 8852 9580
rect 8904 9528 8910 9580
rect 9048 9577 9076 9608
rect 10704 9580 10732 9608
rect 9033 9571 9091 9577
rect 9033 9537 9045 9571
rect 9079 9537 9091 9571
rect 9033 9531 9091 9537
rect 10502 9528 10508 9580
rect 10560 9528 10566 9580
rect 10686 9528 10692 9580
rect 10744 9528 10750 9580
rect 13556 9568 13584 9676
rect 13906 9664 13912 9676
rect 13964 9704 13970 9716
rect 14921 9707 14979 9713
rect 14921 9704 14933 9707
rect 13964 9676 14933 9704
rect 13964 9664 13970 9676
rect 14921 9673 14933 9676
rect 14967 9673 14979 9707
rect 14921 9667 14979 9673
rect 17402 9664 17408 9716
rect 17460 9664 17466 9716
rect 19337 9707 19395 9713
rect 19337 9673 19349 9707
rect 19383 9673 19395 9707
rect 19337 9667 19395 9673
rect 15841 9639 15899 9645
rect 15841 9605 15853 9639
rect 15887 9636 15899 9639
rect 16850 9636 16856 9648
rect 15887 9608 16856 9636
rect 15887 9605 15899 9608
rect 15841 9599 15899 9605
rect 16850 9596 16856 9608
rect 16908 9596 16914 9648
rect 18417 9639 18475 9645
rect 18417 9605 18429 9639
rect 18463 9636 18475 9639
rect 19352 9636 19380 9667
rect 20806 9664 20812 9716
rect 20864 9664 20870 9716
rect 21269 9707 21327 9713
rect 21269 9673 21281 9707
rect 21315 9704 21327 9707
rect 21358 9704 21364 9716
rect 21315 9676 21364 9704
rect 21315 9673 21327 9676
rect 21269 9667 21327 9673
rect 21358 9664 21364 9676
rect 21416 9664 21422 9716
rect 22462 9664 22468 9716
rect 22520 9704 22526 9716
rect 22741 9707 22799 9713
rect 22741 9704 22753 9707
rect 22520 9676 22753 9704
rect 22520 9664 22526 9676
rect 22741 9673 22753 9676
rect 22787 9673 22799 9707
rect 22741 9667 22799 9673
rect 18463 9608 19380 9636
rect 18463 9605 18475 9608
rect 18417 9599 18475 9605
rect 13372 9540 13584 9568
rect 5813 9503 5871 9509
rect 5813 9500 5825 9503
rect 5736 9472 5825 9500
rect 5629 9463 5687 9469
rect 5813 9469 5825 9472
rect 5859 9469 5871 9503
rect 5813 9463 5871 9469
rect 4706 9392 4712 9444
rect 4764 9432 4770 9444
rect 5261 9435 5319 9441
rect 5261 9432 5273 9435
rect 4764 9404 5273 9432
rect 4764 9392 4770 9404
rect 5261 9401 5273 9404
rect 5307 9401 5319 9435
rect 5460 9432 5488 9460
rect 5644 9432 5672 9463
rect 12894 9460 12900 9512
rect 12952 9460 12958 9512
rect 13372 9509 13400 9540
rect 15378 9528 15384 9580
rect 15436 9568 15442 9580
rect 15436 9540 16896 9568
rect 15436 9528 15442 9540
rect 13173 9503 13231 9509
rect 13173 9469 13185 9503
rect 13219 9469 13231 9503
rect 13173 9463 13231 9469
rect 13357 9503 13415 9509
rect 13357 9469 13369 9503
rect 13403 9469 13415 9503
rect 13357 9463 13415 9469
rect 13541 9503 13599 9509
rect 13541 9469 13553 9503
rect 13587 9500 13599 9503
rect 13630 9500 13636 9512
rect 13587 9472 13636 9500
rect 13587 9469 13599 9472
rect 13541 9463 13599 9469
rect 5460 9404 5672 9432
rect 5261 9395 5319 9401
rect 5077 9367 5135 9373
rect 5077 9333 5089 9367
rect 5123 9364 5135 9367
rect 5718 9364 5724 9376
rect 5123 9336 5724 9364
rect 5123 9333 5135 9336
rect 5077 9327 5135 9333
rect 5718 9324 5724 9336
rect 5776 9324 5782 9376
rect 5813 9367 5871 9373
rect 5813 9333 5825 9367
rect 5859 9364 5871 9367
rect 6270 9364 6276 9376
rect 5859 9336 6276 9364
rect 5859 9333 5871 9336
rect 5813 9327 5871 9333
rect 6270 9324 6276 9336
rect 6328 9324 6334 9376
rect 8386 9324 8392 9376
rect 8444 9324 8450 9376
rect 8754 9324 8760 9376
rect 8812 9324 8818 9376
rect 10042 9324 10048 9376
rect 10100 9324 10106 9376
rect 10413 9367 10471 9373
rect 10413 9333 10425 9367
rect 10459 9364 10471 9367
rect 10778 9364 10784 9376
rect 10459 9336 10784 9364
rect 10459 9333 10471 9336
rect 10413 9327 10471 9333
rect 10778 9324 10784 9336
rect 10836 9324 10842 9376
rect 13188 9364 13216 9463
rect 13630 9460 13636 9472
rect 13688 9460 13694 9512
rect 13814 9509 13820 9512
rect 13808 9500 13820 9509
rect 13775 9472 13820 9500
rect 13808 9463 13820 9472
rect 13814 9460 13820 9463
rect 13872 9460 13878 9512
rect 15565 9503 15623 9509
rect 15565 9469 15577 9503
rect 15611 9500 15623 9503
rect 15746 9500 15752 9512
rect 15611 9472 15752 9500
rect 15611 9469 15623 9472
rect 15565 9463 15623 9469
rect 13265 9435 13323 9441
rect 13265 9401 13277 9435
rect 13311 9432 13323 9435
rect 15580 9432 15608 9463
rect 15746 9460 15752 9472
rect 15804 9460 15810 9512
rect 15838 9460 15844 9512
rect 15896 9500 15902 9512
rect 16393 9503 16451 9509
rect 16393 9500 16405 9503
rect 15896 9472 16405 9500
rect 15896 9460 15902 9472
rect 16393 9469 16405 9472
rect 16439 9500 16451 9503
rect 16482 9500 16488 9512
rect 16439 9472 16488 9500
rect 16439 9469 16451 9472
rect 16393 9463 16451 9469
rect 16482 9460 16488 9472
rect 16540 9460 16546 9512
rect 16574 9460 16580 9512
rect 16632 9460 16638 9512
rect 16666 9460 16672 9512
rect 16724 9460 16730 9512
rect 13311 9404 15608 9432
rect 16868 9432 16896 9540
rect 18138 9528 18144 9580
rect 18196 9568 18202 9580
rect 20441 9571 20499 9577
rect 18196 9540 18552 9568
rect 18196 9528 18202 9540
rect 16945 9503 17003 9509
rect 16945 9469 16957 9503
rect 16991 9500 17003 9503
rect 17037 9503 17095 9509
rect 17037 9500 17049 9503
rect 16991 9472 17049 9500
rect 16991 9469 17003 9472
rect 16945 9463 17003 9469
rect 17037 9469 17049 9472
rect 17083 9500 17095 9503
rect 18046 9500 18052 9512
rect 17083 9472 18052 9500
rect 17083 9469 17095 9472
rect 17037 9463 17095 9469
rect 18046 9460 18052 9472
rect 18104 9500 18110 9512
rect 18524 9509 18552 9540
rect 20441 9537 20453 9571
rect 20487 9568 20499 9571
rect 20487 9540 21128 9568
rect 20487 9537 20499 9540
rect 20441 9531 20499 9537
rect 18325 9503 18383 9509
rect 18325 9500 18337 9503
rect 18104 9472 18337 9500
rect 18104 9460 18110 9472
rect 18325 9469 18337 9472
rect 18371 9469 18383 9503
rect 18325 9463 18383 9469
rect 18509 9503 18567 9509
rect 18509 9469 18521 9503
rect 18555 9500 18567 9503
rect 18877 9503 18935 9509
rect 18877 9500 18889 9503
rect 18555 9472 18889 9500
rect 18555 9469 18567 9472
rect 18509 9463 18567 9469
rect 18877 9469 18889 9472
rect 18923 9469 18935 9503
rect 20625 9503 20683 9509
rect 18877 9463 18935 9469
rect 18984 9472 19564 9500
rect 17405 9435 17463 9441
rect 17405 9432 17417 9435
rect 16868 9404 17417 9432
rect 13311 9401 13323 9404
rect 13265 9395 13323 9401
rect 17405 9401 17417 9404
rect 17451 9432 17463 9435
rect 18340 9432 18368 9463
rect 18693 9435 18751 9441
rect 18693 9432 18705 9435
rect 17451 9404 18276 9432
rect 18340 9404 18705 9432
rect 17451 9401 17463 9404
rect 17405 9395 17463 9401
rect 14090 9364 14096 9376
rect 13188 9336 14096 9364
rect 14090 9324 14096 9336
rect 14148 9324 14154 9376
rect 15654 9324 15660 9376
rect 15712 9324 15718 9376
rect 16761 9367 16819 9373
rect 16761 9333 16773 9367
rect 16807 9364 16819 9367
rect 16850 9364 16856 9376
rect 16807 9336 16856 9364
rect 16807 9333 16819 9336
rect 16761 9327 16819 9333
rect 16850 9324 16856 9336
rect 16908 9324 16914 9376
rect 17494 9324 17500 9376
rect 17552 9364 17558 9376
rect 17589 9367 17647 9373
rect 17589 9364 17601 9367
rect 17552 9336 17601 9364
rect 17552 9324 17558 9336
rect 17589 9333 17601 9336
rect 17635 9333 17647 9367
rect 18248 9364 18276 9404
rect 18693 9401 18705 9404
rect 18739 9401 18751 9435
rect 18984 9432 19012 9472
rect 19536 9441 19564 9472
rect 20625 9469 20637 9503
rect 20671 9500 20683 9503
rect 20898 9500 20904 9512
rect 20671 9472 20904 9500
rect 20671 9469 20683 9472
rect 20625 9463 20683 9469
rect 20898 9460 20904 9472
rect 20956 9460 20962 9512
rect 18693 9395 18751 9401
rect 18800 9404 19012 9432
rect 19061 9435 19119 9441
rect 18800 9364 18828 9404
rect 19061 9401 19073 9435
rect 19107 9432 19119 9435
rect 19305 9435 19363 9441
rect 19305 9432 19317 9435
rect 19107 9404 19317 9432
rect 19107 9401 19119 9404
rect 19061 9395 19119 9401
rect 19305 9401 19317 9404
rect 19351 9401 19363 9435
rect 19305 9395 19363 9401
rect 19521 9435 19579 9441
rect 19521 9401 19533 9435
rect 19567 9432 19579 9435
rect 20714 9432 20720 9444
rect 19567 9404 20720 9432
rect 19567 9401 19579 9404
rect 19521 9395 19579 9401
rect 20714 9392 20720 9404
rect 20772 9392 20778 9444
rect 21100 9441 21128 9540
rect 21174 9528 21180 9580
rect 21232 9568 21238 9580
rect 21361 9571 21419 9577
rect 21361 9568 21373 9571
rect 21232 9540 21373 9568
rect 21232 9528 21238 9540
rect 21361 9537 21373 9540
rect 21407 9537 21419 9571
rect 21361 9531 21419 9537
rect 21085 9435 21143 9441
rect 21085 9401 21097 9435
rect 21131 9401 21143 9435
rect 21085 9395 21143 9401
rect 18248 9336 18828 9364
rect 17589 9327 17647 9333
rect 19150 9324 19156 9376
rect 19208 9324 19214 9376
rect 21100 9364 21128 9395
rect 21266 9392 21272 9444
rect 21324 9432 21330 9444
rect 21606 9435 21664 9441
rect 21606 9432 21618 9435
rect 21324 9404 21618 9432
rect 21324 9392 21330 9404
rect 21606 9401 21618 9404
rect 21652 9401 21664 9435
rect 21606 9395 21664 9401
rect 22462 9364 22468 9376
rect 21100 9336 22468 9364
rect 22462 9324 22468 9336
rect 22520 9324 22526 9376
rect 552 9274 23368 9296
rect 552 9222 4322 9274
rect 4374 9222 4386 9274
rect 4438 9222 4450 9274
rect 4502 9222 4514 9274
rect 4566 9222 4578 9274
rect 4630 9222 23368 9274
rect 552 9200 23368 9222
rect 8754 9120 8760 9172
rect 8812 9160 8818 9172
rect 9125 9163 9183 9169
rect 9125 9160 9137 9163
rect 8812 9132 9137 9160
rect 8812 9120 8818 9132
rect 9125 9129 9137 9132
rect 9171 9129 9183 9163
rect 9125 9123 9183 9129
rect 10778 9120 10784 9172
rect 10836 9120 10842 9172
rect 14553 9163 14611 9169
rect 14553 9129 14565 9163
rect 14599 9160 14611 9163
rect 15654 9160 15660 9172
rect 14599 9132 15660 9160
rect 14599 9129 14611 9132
rect 14553 9123 14611 9129
rect 15654 9120 15660 9132
rect 15712 9120 15718 9172
rect 15933 9163 15991 9169
rect 15933 9129 15945 9163
rect 15979 9160 15991 9163
rect 17402 9160 17408 9172
rect 15979 9132 17408 9160
rect 15979 9129 15991 9132
rect 15933 9123 15991 9129
rect 17402 9120 17408 9132
rect 17460 9120 17466 9172
rect 18138 9120 18144 9172
rect 18196 9120 18202 9172
rect 19334 9120 19340 9172
rect 19392 9120 19398 9172
rect 22554 9120 22560 9172
rect 22612 9160 22618 9172
rect 22649 9163 22707 9169
rect 22649 9160 22661 9163
rect 22612 9132 22661 9160
rect 22612 9120 22618 9132
rect 22649 9129 22661 9132
rect 22695 9129 22707 9163
rect 22649 9123 22707 9129
rect 3513 9095 3571 9101
rect 3513 9092 3525 9095
rect 3068 9064 3525 9092
rect 3068 9036 3096 9064
rect 3513 9061 3525 9064
rect 3559 9061 3571 9095
rect 3513 9055 3571 9061
rect 8012 9095 8070 9101
rect 8012 9061 8024 9095
rect 8058 9092 8070 9095
rect 8386 9092 8392 9104
rect 8058 9064 8392 9092
rect 8058 9061 8070 9064
rect 8012 9055 8070 9061
rect 8386 9052 8392 9064
rect 8444 9052 8450 9104
rect 9668 9095 9726 9101
rect 9668 9061 9680 9095
rect 9714 9092 9726 9095
rect 10042 9092 10048 9104
rect 9714 9064 10048 9092
rect 9714 9061 9726 9064
rect 9668 9055 9726 9061
rect 10042 9052 10048 9064
rect 10100 9052 10106 9104
rect 10796 9092 10824 9120
rect 10796 9064 11744 9092
rect 3050 8984 3056 9036
rect 3108 8984 3114 9036
rect 3237 9027 3295 9033
rect 3237 8993 3249 9027
rect 3283 9024 3295 9027
rect 3326 9024 3332 9036
rect 3283 8996 3332 9024
rect 3283 8993 3295 8996
rect 3237 8987 3295 8993
rect 3326 8984 3332 8996
rect 3384 8984 3390 9036
rect 3973 9027 4031 9033
rect 3973 8993 3985 9027
rect 4019 8993 4031 9027
rect 3973 8987 4031 8993
rect 3510 8916 3516 8968
rect 3568 8956 3574 8968
rect 3988 8956 4016 8987
rect 4154 8984 4160 9036
rect 4212 9024 4218 9036
rect 4617 9027 4675 9033
rect 4617 9024 4629 9027
rect 4212 8996 4629 9024
rect 4212 8984 4218 8996
rect 4617 8993 4629 8996
rect 4663 8993 4675 9027
rect 4617 8987 4675 8993
rect 4982 8984 4988 9036
rect 5040 9024 5046 9036
rect 5077 9027 5135 9033
rect 5077 9024 5089 9027
rect 5040 8996 5089 9024
rect 5040 8984 5046 8996
rect 5077 8993 5089 8996
rect 5123 8993 5135 9027
rect 5077 8987 5135 8993
rect 7745 9027 7803 9033
rect 7745 8993 7757 9027
rect 7791 9024 7803 9027
rect 8846 9024 8852 9036
rect 7791 8996 8852 9024
rect 7791 8993 7803 8996
rect 7745 8987 7803 8993
rect 8846 8984 8852 8996
rect 8904 9024 8910 9036
rect 9398 9024 9404 9036
rect 8904 8996 9404 9024
rect 8904 8984 8910 8996
rect 9398 8984 9404 8996
rect 9456 8984 9462 9036
rect 11422 8984 11428 9036
rect 11480 8984 11486 9036
rect 11716 9033 11744 9064
rect 12894 9052 12900 9104
rect 12952 9092 12958 9104
rect 12952 9064 14412 9092
rect 12952 9052 12958 9064
rect 11701 9027 11759 9033
rect 11701 8993 11713 9027
rect 11747 8993 11759 9027
rect 11701 8987 11759 8993
rect 14090 8984 14096 9036
rect 14148 8984 14154 9036
rect 14384 9033 14412 9064
rect 19150 9052 19156 9104
rect 19208 9092 19214 9104
rect 19254 9095 19312 9101
rect 19254 9092 19266 9095
rect 19208 9064 19266 9092
rect 19208 9052 19214 9064
rect 19254 9061 19266 9064
rect 19300 9061 19312 9095
rect 19254 9055 19312 9061
rect 14369 9027 14427 9033
rect 14369 8993 14381 9027
rect 14415 8993 14427 9027
rect 14369 8987 14427 8993
rect 15562 8984 15568 9036
rect 15620 8984 15626 9036
rect 15749 9027 15807 9033
rect 15749 8993 15761 9027
rect 15795 9024 15807 9027
rect 15795 8996 16436 9024
rect 15795 8993 15807 8996
rect 15749 8987 15807 8993
rect 3568 8928 4016 8956
rect 3568 8916 3574 8928
rect 4062 8916 4068 8968
rect 4120 8916 4126 8968
rect 4893 8959 4951 8965
rect 4893 8956 4905 8959
rect 4356 8928 4905 8956
rect 4356 8897 4384 8928
rect 4893 8925 4905 8928
rect 4939 8925 4951 8959
rect 4893 8919 4951 8925
rect 11238 8916 11244 8968
rect 11296 8956 11302 8968
rect 11517 8959 11575 8965
rect 11517 8956 11529 8959
rect 11296 8928 11529 8956
rect 11296 8916 11302 8928
rect 11517 8925 11529 8928
rect 11563 8956 11575 8959
rect 11606 8956 11612 8968
rect 11563 8928 11612 8956
rect 11563 8925 11575 8928
rect 11517 8919 11575 8925
rect 11606 8916 11612 8928
rect 11664 8916 11670 8968
rect 13906 8916 13912 8968
rect 13964 8956 13970 8968
rect 14185 8959 14243 8965
rect 14185 8956 14197 8959
rect 13964 8928 14197 8956
rect 13964 8916 13970 8928
rect 14185 8925 14197 8928
rect 14231 8925 14243 8959
rect 14185 8919 14243 8925
rect 4341 8891 4399 8897
rect 4341 8857 4353 8891
rect 4387 8857 4399 8891
rect 4341 8851 4399 8857
rect 13814 8848 13820 8900
rect 13872 8888 13878 8900
rect 13998 8888 14004 8900
rect 13872 8860 14004 8888
rect 13872 8848 13878 8860
rect 13998 8848 14004 8860
rect 14056 8888 14062 8900
rect 15746 8888 15752 8900
rect 14056 8860 15752 8888
rect 14056 8848 14062 8860
rect 15746 8848 15752 8860
rect 15804 8848 15810 8900
rect 16408 8897 16436 8996
rect 17494 8984 17500 9036
rect 17552 9033 17558 9036
rect 17552 9024 17564 9033
rect 19352 9024 19380 9120
rect 19521 9027 19579 9033
rect 19521 9024 19533 9027
rect 17552 8996 17597 9024
rect 19352 8996 19533 9024
rect 17552 8987 17564 8996
rect 19521 8993 19533 8996
rect 19567 8993 19579 9027
rect 19521 8987 19579 8993
rect 17552 8984 17558 8987
rect 21358 8984 21364 9036
rect 21416 9024 21422 9036
rect 21525 9027 21583 9033
rect 21525 9024 21537 9027
rect 21416 8996 21537 9024
rect 21416 8984 21422 8996
rect 21525 8993 21537 8996
rect 21571 8993 21583 9027
rect 21525 8987 21583 8993
rect 17773 8959 17831 8965
rect 17773 8925 17785 8959
rect 17819 8956 17831 8959
rect 17819 8928 17908 8956
rect 17819 8925 17831 8928
rect 17773 8919 17831 8925
rect 16393 8891 16451 8897
rect 16393 8857 16405 8891
rect 16439 8888 16451 8891
rect 16666 8888 16672 8900
rect 16439 8860 16672 8888
rect 16439 8857 16451 8860
rect 16393 8851 16451 8857
rect 16666 8848 16672 8860
rect 16724 8848 16730 8900
rect 3142 8780 3148 8832
rect 3200 8780 3206 8832
rect 3697 8823 3755 8829
rect 3697 8789 3709 8823
rect 3743 8820 3755 8823
rect 4062 8820 4068 8832
rect 3743 8792 4068 8820
rect 3743 8789 3755 8792
rect 3697 8783 3755 8789
rect 4062 8780 4068 8792
rect 4120 8780 4126 8832
rect 5074 8780 5080 8832
rect 5132 8780 5138 8832
rect 5261 8823 5319 8829
rect 5261 8789 5273 8823
rect 5307 8820 5319 8823
rect 5902 8820 5908 8832
rect 5307 8792 5908 8820
rect 5307 8789 5319 8792
rect 5261 8783 5319 8789
rect 5902 8780 5908 8792
rect 5960 8780 5966 8832
rect 10962 8780 10968 8832
rect 11020 8820 11026 8832
rect 11425 8823 11483 8829
rect 11425 8820 11437 8823
rect 11020 8792 11437 8820
rect 11020 8780 11026 8792
rect 11425 8789 11437 8792
rect 11471 8789 11483 8823
rect 11425 8783 11483 8789
rect 11885 8823 11943 8829
rect 11885 8789 11897 8823
rect 11931 8820 11943 8823
rect 12526 8820 12532 8832
rect 11931 8792 12532 8820
rect 11931 8789 11943 8792
rect 11885 8783 11943 8789
rect 12526 8780 12532 8792
rect 12584 8780 12590 8832
rect 14182 8780 14188 8832
rect 14240 8780 14246 8832
rect 17880 8820 17908 8928
rect 20806 8916 20812 8968
rect 20864 8956 20870 8968
rect 21269 8959 21327 8965
rect 21269 8956 21281 8959
rect 20864 8928 21281 8956
rect 20864 8916 20870 8928
rect 21269 8925 21281 8928
rect 21315 8925 21327 8959
rect 21269 8919 21327 8925
rect 20806 8820 20812 8832
rect 17880 8792 20812 8820
rect 20806 8780 20812 8792
rect 20864 8780 20870 8832
rect 552 8730 23368 8752
rect 552 8678 3662 8730
rect 3714 8678 3726 8730
rect 3778 8678 3790 8730
rect 3842 8678 3854 8730
rect 3906 8678 3918 8730
rect 3970 8678 23368 8730
rect 552 8656 23368 8678
rect 3881 8619 3939 8625
rect 3881 8585 3893 8619
rect 3927 8616 3939 8619
rect 4062 8616 4068 8628
rect 3927 8588 4068 8616
rect 3927 8585 3939 8588
rect 3881 8579 3939 8585
rect 4062 8576 4068 8588
rect 4120 8576 4126 8628
rect 4801 8619 4859 8625
rect 4801 8585 4813 8619
rect 4847 8585 4859 8619
rect 4801 8579 4859 8585
rect 4816 8548 4844 8579
rect 4982 8576 4988 8628
rect 5040 8576 5046 8628
rect 5718 8576 5724 8628
rect 5776 8616 5782 8628
rect 5997 8619 6055 8625
rect 5997 8616 6009 8619
rect 5776 8588 6009 8616
rect 5776 8576 5782 8588
rect 5997 8585 6009 8588
rect 6043 8616 6055 8619
rect 6362 8616 6368 8628
rect 6043 8588 6368 8616
rect 6043 8585 6055 8588
rect 5997 8579 6055 8585
rect 6362 8576 6368 8588
rect 6420 8616 6426 8628
rect 7469 8619 7527 8625
rect 7469 8616 7481 8619
rect 6420 8588 7481 8616
rect 6420 8576 6426 8588
rect 7469 8585 7481 8588
rect 7515 8585 7527 8619
rect 7469 8579 7527 8585
rect 5442 8548 5448 8560
rect 4816 8520 5448 8548
rect 5442 8508 5448 8520
rect 5500 8508 5506 8560
rect 6086 8508 6092 8560
rect 6144 8548 6150 8560
rect 6549 8551 6607 8557
rect 6549 8548 6561 8551
rect 6144 8520 6561 8548
rect 6144 8508 6150 8520
rect 6549 8517 6561 8520
rect 6595 8517 6607 8551
rect 6549 8511 6607 8517
rect 5828 8452 6592 8480
rect 3142 8372 3148 8424
rect 3200 8412 3206 8424
rect 3200 8387 3940 8412
rect 3200 8384 3985 8387
rect 3200 8372 3206 8384
rect 3912 8381 3985 8384
rect 3418 8304 3424 8356
rect 3476 8344 3482 8356
rect 3697 8347 3755 8353
rect 3912 8350 3939 8381
rect 3697 8344 3709 8347
rect 3476 8316 3709 8344
rect 3476 8304 3482 8316
rect 3697 8313 3709 8316
rect 3743 8313 3755 8347
rect 3927 8347 3939 8350
rect 3973 8347 3985 8381
rect 5828 8356 5856 8452
rect 6270 8372 6276 8424
rect 6328 8372 6334 8424
rect 6362 8372 6368 8424
rect 6420 8372 6426 8424
rect 6564 8421 6592 8452
rect 6549 8415 6607 8421
rect 6549 8381 6561 8415
rect 6595 8381 6607 8415
rect 6549 8375 6607 8381
rect 6730 8372 6736 8424
rect 6788 8412 6794 8424
rect 7377 8415 7435 8421
rect 7377 8412 7389 8415
rect 6788 8384 7389 8412
rect 6788 8372 6794 8384
rect 7377 8381 7389 8384
rect 7423 8381 7435 8415
rect 7484 8412 7512 8579
rect 7742 8576 7748 8628
rect 7800 8616 7806 8628
rect 8389 8619 8447 8625
rect 8389 8616 8401 8619
rect 7800 8588 8401 8616
rect 7800 8576 7806 8588
rect 8389 8585 8401 8588
rect 8435 8585 8447 8619
rect 8389 8579 8447 8585
rect 10962 8576 10968 8628
rect 11020 8616 11026 8628
rect 11287 8619 11345 8625
rect 11287 8616 11299 8619
rect 11020 8588 11299 8616
rect 11020 8576 11026 8588
rect 11287 8585 11299 8588
rect 11333 8585 11345 8619
rect 11287 8579 11345 8585
rect 15470 8576 15476 8628
rect 15528 8576 15534 8628
rect 16666 8576 16672 8628
rect 16724 8616 16730 8628
rect 17129 8619 17187 8625
rect 17129 8616 17141 8619
rect 16724 8588 17141 8616
rect 16724 8576 16730 8588
rect 17129 8585 17141 8588
rect 17175 8585 17187 8619
rect 17129 8579 17187 8585
rect 21269 8619 21327 8625
rect 21269 8585 21281 8619
rect 21315 8616 21327 8619
rect 21358 8616 21364 8628
rect 21315 8588 21364 8616
rect 21315 8585 21327 8588
rect 21269 8579 21327 8585
rect 21358 8576 21364 8588
rect 21416 8576 21422 8628
rect 21453 8619 21511 8625
rect 21453 8585 21465 8619
rect 21499 8616 21511 8619
rect 22002 8616 22008 8628
rect 21499 8588 22008 8616
rect 21499 8585 21511 8588
rect 21453 8579 21511 8585
rect 22002 8576 22008 8588
rect 22060 8576 22066 8628
rect 7653 8483 7711 8489
rect 7653 8449 7665 8483
rect 7699 8480 7711 8483
rect 7760 8480 7788 8576
rect 10597 8551 10655 8557
rect 10597 8517 10609 8551
rect 10643 8548 10655 8551
rect 11146 8548 11152 8560
rect 10643 8520 11152 8548
rect 10643 8517 10655 8520
rect 10597 8511 10655 8517
rect 11146 8508 11152 8520
rect 11204 8508 11210 8560
rect 15657 8551 15715 8557
rect 13188 8520 14596 8548
rect 8573 8483 8631 8489
rect 7699 8452 7788 8480
rect 7852 8452 8448 8480
rect 7699 8449 7711 8452
rect 7653 8443 7711 8449
rect 7745 8415 7803 8421
rect 7745 8412 7757 8415
rect 7484 8384 7757 8412
rect 7377 8375 7435 8381
rect 7745 8381 7757 8384
rect 7791 8412 7803 8415
rect 7852 8412 7880 8452
rect 7791 8384 7880 8412
rect 7929 8415 7987 8421
rect 7791 8381 7803 8384
rect 7745 8375 7803 8381
rect 7929 8381 7941 8415
rect 7975 8412 7987 8415
rect 7975 8384 8340 8412
rect 7975 8381 7987 8384
rect 7929 8375 7987 8381
rect 3927 8341 3985 8347
rect 4154 8344 4160 8356
rect 3697 8307 3755 8313
rect 4080 8316 4160 8344
rect 4080 8285 4108 8316
rect 4154 8304 4160 8316
rect 4212 8304 4218 8356
rect 4617 8347 4675 8353
rect 4617 8313 4629 8347
rect 4663 8344 4675 8347
rect 4706 8344 4712 8356
rect 4663 8316 4712 8344
rect 4663 8313 4675 8316
rect 4617 8307 4675 8313
rect 4706 8304 4712 8316
rect 4764 8304 4770 8356
rect 4798 8304 4804 8356
rect 4856 8353 4862 8356
rect 4856 8347 4875 8353
rect 4863 8313 4875 8347
rect 4856 8307 4875 8313
rect 4856 8304 4862 8307
rect 5810 8304 5816 8356
rect 5868 8304 5874 8356
rect 6029 8347 6087 8353
rect 6029 8313 6041 8347
rect 6075 8344 6087 8347
rect 6288 8344 6316 8372
rect 6075 8316 6316 8344
rect 7392 8344 7420 8375
rect 7944 8344 7972 8375
rect 7392 8316 7972 8344
rect 6075 8313 6087 8316
rect 6029 8307 6087 8313
rect 4065 8279 4123 8285
rect 4065 8245 4077 8279
rect 4111 8245 4123 8279
rect 4065 8239 4123 8245
rect 6178 8236 6184 8288
rect 6236 8236 6242 8288
rect 7653 8279 7711 8285
rect 7653 8245 7665 8279
rect 7699 8276 7711 8279
rect 7742 8276 7748 8288
rect 7699 8248 7748 8276
rect 7699 8245 7711 8248
rect 7653 8239 7711 8245
rect 7742 8236 7748 8248
rect 7800 8236 7806 8288
rect 8113 8279 8171 8285
rect 8113 8245 8125 8279
rect 8159 8276 8171 8279
rect 8202 8276 8208 8288
rect 8159 8248 8208 8276
rect 8159 8245 8171 8248
rect 8113 8239 8171 8245
rect 8202 8236 8208 8248
rect 8260 8236 8266 8288
rect 8312 8276 8340 8384
rect 8420 8353 8448 8452
rect 8573 8449 8585 8483
rect 8619 8480 8631 8483
rect 8754 8480 8760 8492
rect 8619 8452 8760 8480
rect 8619 8449 8631 8452
rect 8573 8443 8631 8449
rect 8754 8440 8760 8452
rect 8812 8440 8818 8492
rect 10689 8483 10747 8489
rect 10689 8480 10701 8483
rect 10428 8452 10701 8480
rect 10428 8421 10456 8452
rect 10689 8449 10701 8452
rect 10735 8480 10747 8483
rect 10778 8480 10784 8492
rect 10735 8452 10784 8480
rect 10735 8449 10747 8452
rect 10689 8443 10747 8449
rect 10778 8440 10784 8452
rect 10836 8480 10842 8492
rect 11517 8483 11575 8489
rect 10836 8452 11192 8480
rect 10836 8440 10842 8452
rect 11164 8421 11192 8452
rect 11517 8449 11529 8483
rect 11563 8480 11575 8483
rect 11563 8452 12388 8480
rect 11563 8449 11575 8452
rect 11517 8443 11575 8449
rect 8665 8415 8723 8421
rect 8665 8381 8677 8415
rect 8711 8381 8723 8415
rect 8665 8375 8723 8381
rect 10413 8415 10471 8421
rect 10413 8381 10425 8415
rect 10459 8381 10471 8415
rect 10413 8375 10471 8381
rect 10597 8415 10655 8421
rect 10597 8381 10609 8415
rect 10643 8412 10655 8415
rect 10873 8415 10931 8421
rect 10873 8412 10885 8415
rect 10643 8384 10885 8412
rect 10643 8381 10655 8384
rect 10597 8375 10655 8381
rect 10873 8381 10885 8384
rect 10919 8381 10931 8415
rect 10873 8375 10931 8381
rect 11149 8415 11207 8421
rect 11149 8381 11161 8415
rect 11195 8381 11207 8415
rect 11149 8375 11207 8381
rect 8389 8347 8448 8353
rect 8389 8313 8401 8347
rect 8435 8316 8448 8347
rect 8680 8344 8708 8375
rect 10612 8344 10640 8375
rect 8496 8316 8708 8344
rect 8864 8316 10640 8344
rect 10888 8344 10916 8375
rect 11422 8372 11428 8424
rect 11480 8372 11486 8424
rect 11606 8372 11612 8424
rect 11664 8372 11670 8424
rect 12360 8421 12388 8452
rect 12345 8415 12403 8421
rect 12345 8381 12357 8415
rect 12391 8381 12403 8415
rect 12345 8375 12403 8381
rect 12526 8372 12532 8424
rect 12584 8372 12590 8424
rect 12894 8372 12900 8424
rect 12952 8412 12958 8424
rect 13188 8421 13216 8520
rect 13265 8483 13323 8489
rect 13265 8449 13277 8483
rect 13311 8480 13323 8483
rect 13538 8480 13544 8492
rect 13311 8452 13544 8480
rect 13311 8449 13323 8452
rect 13265 8443 13323 8449
rect 13538 8440 13544 8452
rect 13596 8480 13602 8492
rect 13633 8483 13691 8489
rect 13633 8480 13645 8483
rect 13596 8452 13645 8480
rect 13596 8440 13602 8452
rect 13633 8449 13645 8452
rect 13679 8449 13691 8483
rect 14182 8480 14188 8492
rect 13633 8443 13691 8449
rect 13740 8452 14188 8480
rect 13740 8421 13768 8452
rect 14182 8440 14188 8452
rect 14240 8440 14246 8492
rect 14568 8489 14596 8520
rect 15657 8517 15669 8551
rect 15703 8517 15715 8551
rect 15657 8511 15715 8517
rect 21821 8551 21879 8557
rect 21821 8517 21833 8551
rect 21867 8548 21879 8551
rect 21910 8548 21916 8560
rect 21867 8520 21916 8548
rect 21867 8517 21879 8520
rect 21821 8511 21879 8517
rect 14553 8483 14611 8489
rect 14553 8449 14565 8483
rect 14599 8449 14611 8483
rect 15672 8480 15700 8511
rect 21910 8508 21916 8520
rect 21968 8508 21974 8560
rect 15672 8452 15884 8480
rect 14553 8443 14611 8449
rect 13173 8415 13231 8421
rect 13173 8412 13185 8415
rect 12952 8384 13185 8412
rect 12952 8372 12958 8384
rect 13173 8381 13185 8384
rect 13219 8381 13231 8415
rect 13173 8375 13231 8381
rect 13357 8415 13415 8421
rect 13357 8381 13369 8415
rect 13403 8381 13415 8415
rect 13357 8375 13415 8381
rect 13725 8415 13783 8421
rect 13725 8381 13737 8415
rect 13771 8381 13783 8415
rect 14090 8412 14096 8424
rect 13725 8375 13783 8381
rect 13832 8384 14096 8412
rect 11440 8344 11468 8372
rect 10888 8316 11468 8344
rect 12544 8344 12572 8372
rect 13372 8344 13400 8375
rect 13832 8344 13860 8384
rect 14090 8372 14096 8384
rect 14148 8412 14154 8424
rect 14369 8415 14427 8421
rect 14369 8412 14381 8415
rect 14148 8384 14381 8412
rect 14148 8372 14154 8384
rect 14369 8381 14381 8384
rect 14415 8381 14427 8415
rect 14369 8375 14427 8381
rect 15105 8415 15163 8421
rect 15105 8381 15117 8415
rect 15151 8381 15163 8415
rect 15105 8375 15163 8381
rect 12544 8316 13860 8344
rect 8435 8313 8447 8316
rect 8389 8307 8447 8313
rect 8496 8276 8524 8316
rect 8864 8285 8892 8316
rect 14182 8304 14188 8356
rect 14240 8304 14246 8356
rect 15120 8344 15148 8375
rect 15746 8372 15752 8424
rect 15804 8372 15810 8424
rect 15856 8412 15884 8452
rect 16005 8415 16063 8421
rect 16005 8412 16017 8415
rect 15856 8384 16017 8412
rect 16005 8381 16017 8384
rect 16051 8381 16063 8415
rect 16005 8375 16063 8381
rect 15562 8344 15568 8356
rect 15120 8316 15568 8344
rect 15562 8304 15568 8316
rect 15620 8344 15626 8356
rect 16206 8344 16212 8356
rect 15620 8316 16212 8344
rect 15620 8304 15626 8316
rect 16206 8304 16212 8316
rect 16264 8304 16270 8356
rect 20990 8304 20996 8356
rect 21048 8344 21054 8356
rect 21266 8344 21272 8356
rect 21048 8316 21272 8344
rect 21048 8304 21054 8316
rect 21266 8304 21272 8316
rect 21324 8344 21330 8356
rect 21453 8347 21511 8353
rect 21453 8344 21465 8347
rect 21324 8316 21465 8344
rect 21324 8304 21330 8316
rect 21453 8313 21465 8316
rect 21499 8313 21511 8347
rect 21453 8307 21511 8313
rect 8312 8248 8524 8276
rect 8849 8279 8907 8285
rect 8849 8245 8861 8279
rect 8895 8245 8907 8279
rect 8849 8239 8907 8245
rect 11057 8279 11115 8285
rect 11057 8245 11069 8279
rect 11103 8276 11115 8279
rect 11606 8276 11612 8288
rect 11103 8248 11612 8276
rect 11103 8245 11115 8248
rect 11057 8239 11115 8245
rect 11606 8236 11612 8248
rect 11664 8236 11670 8288
rect 12529 8279 12587 8285
rect 12529 8245 12541 8279
rect 12575 8276 12587 8279
rect 12802 8276 12808 8288
rect 12575 8248 12808 8276
rect 12575 8245 12587 8248
rect 12529 8239 12587 8245
rect 12802 8236 12808 8248
rect 12860 8236 12866 8288
rect 14093 8279 14151 8285
rect 14093 8245 14105 8279
rect 14139 8276 14151 8279
rect 14458 8276 14464 8288
rect 14139 8248 14464 8276
rect 14139 8245 14151 8248
rect 14093 8239 14151 8245
rect 14458 8236 14464 8248
rect 14516 8236 14522 8288
rect 15378 8236 15384 8288
rect 15436 8276 15442 8288
rect 15473 8279 15531 8285
rect 15473 8276 15485 8279
rect 15436 8248 15485 8276
rect 15436 8236 15442 8248
rect 15473 8245 15485 8248
rect 15519 8245 15531 8279
rect 15473 8239 15531 8245
rect 19150 8236 19156 8288
rect 19208 8276 19214 8288
rect 21008 8276 21036 8304
rect 19208 8248 21036 8276
rect 19208 8236 19214 8248
rect 552 8186 23368 8208
rect 552 8134 4322 8186
rect 4374 8134 4386 8186
rect 4438 8134 4450 8186
rect 4502 8134 4514 8186
rect 4566 8134 4578 8186
rect 4630 8134 23368 8186
rect 552 8112 23368 8134
rect 3142 8032 3148 8084
rect 3200 8072 3206 8084
rect 3510 8072 3516 8084
rect 3200 8044 3516 8072
rect 3200 8032 3206 8044
rect 3510 8032 3516 8044
rect 3568 8072 3574 8084
rect 3973 8075 4031 8081
rect 3973 8072 3985 8075
rect 3568 8044 3985 8072
rect 3568 8032 3574 8044
rect 3973 8041 3985 8044
rect 4019 8041 4031 8075
rect 3973 8035 4031 8041
rect 4065 8075 4123 8081
rect 4065 8041 4077 8075
rect 4111 8072 4123 8075
rect 4706 8072 4712 8084
rect 4111 8044 4712 8072
rect 4111 8041 4123 8044
rect 4065 8035 4123 8041
rect 4706 8032 4712 8044
rect 4764 8032 4770 8084
rect 6273 8075 6331 8081
rect 6273 8041 6285 8075
rect 6319 8072 6331 8075
rect 6319 8044 6914 8072
rect 6319 8041 6331 8044
rect 6273 8035 6331 8041
rect 2685 8007 2743 8013
rect 2685 7973 2697 8007
rect 2731 8004 2743 8007
rect 3050 8004 3056 8016
rect 2731 7976 3056 8004
rect 2731 7973 2743 7976
rect 2685 7967 2743 7973
rect 2225 7939 2283 7945
rect 2225 7905 2237 7939
rect 2271 7905 2283 7939
rect 2225 7899 2283 7905
rect 2409 7939 2467 7945
rect 2409 7905 2421 7939
rect 2455 7936 2467 7939
rect 2700 7936 2728 7967
rect 3050 7964 3056 7976
rect 3108 8004 3114 8016
rect 3789 8007 3847 8013
rect 3789 8004 3801 8007
rect 3108 7976 3801 8004
rect 3108 7964 3114 7976
rect 3344 7948 3372 7976
rect 3789 7973 3801 7976
rect 3835 7973 3847 8007
rect 6886 8004 6914 8044
rect 15470 8032 15476 8084
rect 15528 8072 15534 8084
rect 16117 8075 16175 8081
rect 16117 8072 16129 8075
rect 15528 8044 16129 8072
rect 15528 8032 15534 8044
rect 16117 8041 16129 8044
rect 16163 8041 16175 8075
rect 16117 8035 16175 8041
rect 16206 8032 16212 8084
rect 16264 8072 16270 8084
rect 16850 8081 16856 8084
rect 16669 8075 16727 8081
rect 16669 8072 16681 8075
rect 16264 8044 16681 8072
rect 16264 8032 16270 8044
rect 16669 8041 16681 8044
rect 16715 8041 16727 8075
rect 16669 8035 16727 8041
rect 16837 8075 16856 8081
rect 16837 8041 16849 8075
rect 16837 8035 16856 8041
rect 16850 8032 16856 8035
rect 16908 8032 16914 8084
rect 21269 8075 21327 8081
rect 21269 8041 21281 8075
rect 21315 8072 21327 8075
rect 21450 8072 21456 8084
rect 21315 8044 21456 8072
rect 21315 8041 21327 8044
rect 21269 8035 21327 8041
rect 21450 8032 21456 8044
rect 21508 8032 21514 8084
rect 7837 8007 7895 8013
rect 7837 8004 7849 8007
rect 6886 7976 7849 8004
rect 3789 7967 3847 7973
rect 7837 7973 7849 7976
rect 7883 7973 7895 8007
rect 14182 8004 14188 8016
rect 7837 7967 7895 7973
rect 13740 7976 14188 8004
rect 2455 7908 2728 7936
rect 2869 7939 2927 7945
rect 2455 7905 2467 7908
rect 2409 7899 2467 7905
rect 2869 7905 2881 7939
rect 2915 7905 2927 7939
rect 2869 7899 2927 7905
rect 2240 7868 2268 7899
rect 2884 7868 2912 7899
rect 3142 7896 3148 7948
rect 3200 7896 3206 7948
rect 3326 7896 3332 7948
rect 3384 7896 3390 7948
rect 3418 7896 3424 7948
rect 3476 7896 3482 7948
rect 4157 7939 4215 7945
rect 4157 7905 4169 7939
rect 4203 7905 4215 7939
rect 4157 7899 4215 7905
rect 3436 7868 3464 7896
rect 4172 7868 4200 7899
rect 5902 7896 5908 7948
rect 5960 7896 5966 7948
rect 6089 7939 6147 7945
rect 6089 7905 6101 7939
rect 6135 7936 6147 7939
rect 6178 7936 6184 7948
rect 6135 7908 6184 7936
rect 6135 7905 6147 7908
rect 6089 7899 6147 7905
rect 6178 7896 6184 7908
rect 6236 7896 6242 7948
rect 6549 7939 6607 7945
rect 6549 7905 6561 7939
rect 6595 7936 6607 7939
rect 6730 7936 6736 7948
rect 6595 7908 6736 7936
rect 6595 7905 6607 7908
rect 6549 7899 6607 7905
rect 6730 7896 6736 7908
rect 6788 7896 6794 7948
rect 8113 7939 8171 7945
rect 8113 7905 8125 7939
rect 8159 7936 8171 7939
rect 8386 7936 8392 7948
rect 8159 7908 8392 7936
rect 8159 7905 8171 7908
rect 8113 7899 8171 7905
rect 8386 7896 8392 7908
rect 8444 7896 8450 7948
rect 8573 7939 8631 7945
rect 8573 7905 8585 7939
rect 8619 7936 8631 7939
rect 8754 7936 8760 7948
rect 8619 7908 8760 7936
rect 8619 7905 8631 7908
rect 8573 7899 8631 7905
rect 8754 7896 8760 7908
rect 8812 7896 8818 7948
rect 10962 7896 10968 7948
rect 11020 7936 11026 7948
rect 11333 7939 11391 7945
rect 11333 7936 11345 7939
rect 11020 7908 11345 7936
rect 11020 7896 11026 7908
rect 11333 7905 11345 7908
rect 11379 7905 11391 7939
rect 11333 7899 11391 7905
rect 11606 7896 11612 7948
rect 11664 7896 11670 7948
rect 11793 7939 11851 7945
rect 11793 7905 11805 7939
rect 11839 7905 11851 7939
rect 11793 7899 11851 7905
rect 2240 7840 4200 7868
rect 6362 7828 6368 7880
rect 6420 7868 6426 7880
rect 6457 7871 6515 7877
rect 6457 7868 6469 7871
rect 6420 7840 6469 7868
rect 6420 7828 6426 7840
rect 6457 7837 6469 7840
rect 6503 7837 6515 7871
rect 6457 7831 6515 7837
rect 7374 7828 7380 7880
rect 7432 7868 7438 7880
rect 7929 7871 7987 7877
rect 7929 7868 7941 7871
rect 7432 7840 7941 7868
rect 7432 7828 7438 7840
rect 7929 7837 7941 7840
rect 7975 7837 7987 7871
rect 7929 7831 7987 7837
rect 8202 7828 8208 7880
rect 8260 7868 8266 7880
rect 8481 7871 8539 7877
rect 8481 7868 8493 7871
rect 8260 7840 8493 7868
rect 8260 7828 8266 7840
rect 8481 7837 8493 7840
rect 8527 7837 8539 7871
rect 8481 7831 8539 7837
rect 11146 7828 11152 7880
rect 11204 7868 11210 7880
rect 11241 7871 11299 7877
rect 11241 7868 11253 7871
rect 11204 7840 11253 7868
rect 11204 7828 11210 7840
rect 11241 7837 11253 7840
rect 11287 7868 11299 7871
rect 11808 7868 11836 7899
rect 13538 7896 13544 7948
rect 13596 7896 13602 7948
rect 13740 7945 13768 7976
rect 14182 7964 14188 7976
rect 14240 7964 14246 8016
rect 16482 7964 16488 8016
rect 16540 8004 16546 8016
rect 17037 8007 17095 8013
rect 17037 8004 17049 8007
rect 16540 7976 17049 8004
rect 16540 7964 16546 7976
rect 17037 7973 17049 7976
rect 17083 7973 17095 8007
rect 19242 8004 19248 8016
rect 17037 7967 17095 7973
rect 18708 7976 19248 8004
rect 13725 7939 13783 7945
rect 13725 7905 13737 7939
rect 13771 7905 13783 7939
rect 13725 7899 13783 7905
rect 13906 7896 13912 7948
rect 13964 7936 13970 7948
rect 14001 7939 14059 7945
rect 14001 7936 14013 7939
rect 13964 7908 14013 7936
rect 13964 7896 13970 7908
rect 14001 7905 14013 7908
rect 14047 7905 14059 7939
rect 14001 7899 14059 7905
rect 14274 7896 14280 7948
rect 14332 7896 14338 7948
rect 16301 7939 16359 7945
rect 16301 7905 16313 7939
rect 16347 7905 16359 7939
rect 16301 7899 16359 7905
rect 16577 7939 16635 7945
rect 16577 7905 16589 7939
rect 16623 7936 16635 7939
rect 16850 7936 16856 7948
rect 16623 7908 16856 7936
rect 16623 7905 16635 7908
rect 16577 7899 16635 7905
rect 11287 7840 11836 7868
rect 11287 7837 11299 7840
rect 11241 7831 11299 7837
rect 13262 7828 13268 7880
rect 13320 7868 13326 7880
rect 14093 7871 14151 7877
rect 14093 7868 14105 7871
rect 13320 7840 14105 7868
rect 13320 7828 13326 7840
rect 14093 7837 14105 7840
rect 14139 7837 14151 7871
rect 16316 7868 16344 7899
rect 16850 7896 16856 7908
rect 16908 7896 16914 7948
rect 18322 7896 18328 7948
rect 18380 7936 18386 7948
rect 18708 7945 18736 7976
rect 19242 7964 19248 7976
rect 19300 7964 19306 8016
rect 21818 8004 21824 8016
rect 21652 7976 21824 8004
rect 18693 7939 18751 7945
rect 18693 7936 18705 7939
rect 18380 7908 18705 7936
rect 18380 7896 18386 7908
rect 18693 7905 18705 7908
rect 18739 7905 18751 7939
rect 18693 7899 18751 7905
rect 18782 7896 18788 7948
rect 18840 7936 18846 7948
rect 21652 7945 21680 7976
rect 21818 7964 21824 7976
rect 21876 8004 21882 8016
rect 22097 8007 22155 8013
rect 22097 8004 22109 8007
rect 21876 7976 22109 8004
rect 21876 7964 21882 7976
rect 22097 7973 22109 7976
rect 22143 7973 22155 8007
rect 22097 7967 22155 7973
rect 18949 7939 19007 7945
rect 18949 7936 18961 7939
rect 18840 7908 18961 7936
rect 18840 7896 18846 7908
rect 18949 7905 18961 7908
rect 18995 7905 19007 7939
rect 18949 7899 19007 7905
rect 21637 7939 21695 7945
rect 21637 7905 21649 7939
rect 21683 7905 21695 7939
rect 21637 7899 21695 7905
rect 21910 7896 21916 7948
rect 21968 7896 21974 7948
rect 16666 7868 16672 7880
rect 16316 7840 16672 7868
rect 14093 7831 14151 7837
rect 16666 7828 16672 7840
rect 16724 7828 16730 7880
rect 21450 7828 21456 7880
rect 21508 7828 21514 7880
rect 21545 7871 21603 7877
rect 21545 7837 21557 7871
rect 21591 7837 21603 7871
rect 21545 7831 21603 7837
rect 21729 7871 21787 7877
rect 21729 7837 21741 7871
rect 21775 7868 21787 7871
rect 22830 7868 22836 7880
rect 21775 7840 22836 7868
rect 21775 7837 21787 7840
rect 21729 7831 21787 7837
rect 8941 7803 8999 7809
rect 8941 7769 8953 7803
rect 8987 7800 8999 7803
rect 9490 7800 9496 7812
rect 8987 7772 9496 7800
rect 8987 7769 8999 7772
rect 8941 7763 8999 7769
rect 9490 7760 9496 7772
rect 9548 7760 9554 7812
rect 2314 7692 2320 7744
rect 2372 7692 2378 7744
rect 2406 7692 2412 7744
rect 2464 7732 2470 7744
rect 2501 7735 2559 7741
rect 2501 7732 2513 7735
rect 2464 7704 2513 7732
rect 2464 7692 2470 7704
rect 2501 7701 2513 7704
rect 2547 7701 2559 7735
rect 2501 7695 2559 7701
rect 2958 7692 2964 7744
rect 3016 7692 3022 7744
rect 4246 7692 4252 7744
rect 4304 7732 4310 7744
rect 4341 7735 4399 7741
rect 4341 7732 4353 7735
rect 4304 7704 4353 7732
rect 4304 7692 4310 7704
rect 4341 7701 4353 7704
rect 4387 7701 4399 7735
rect 4341 7695 4399 7701
rect 6086 7692 6092 7744
rect 6144 7692 6150 7744
rect 6914 7692 6920 7744
rect 6972 7692 6978 7744
rect 7926 7692 7932 7744
rect 7984 7692 7990 7744
rect 8297 7735 8355 7741
rect 8297 7701 8309 7735
rect 8343 7732 8355 7735
rect 9766 7732 9772 7744
rect 8343 7704 9772 7732
rect 8343 7701 8355 7704
rect 8297 7695 8355 7701
rect 9766 7692 9772 7704
rect 9824 7692 9830 7744
rect 11054 7692 11060 7744
rect 11112 7692 11118 7744
rect 11606 7692 11612 7744
rect 11664 7692 11670 7744
rect 13630 7692 13636 7744
rect 13688 7732 13694 7744
rect 13725 7735 13783 7741
rect 13725 7732 13737 7735
rect 13688 7704 13737 7732
rect 13688 7692 13694 7704
rect 13725 7701 13737 7704
rect 13771 7701 13783 7735
rect 13725 7695 13783 7701
rect 13998 7692 14004 7744
rect 14056 7692 14062 7744
rect 14461 7735 14519 7741
rect 14461 7701 14473 7735
rect 14507 7732 14519 7735
rect 16574 7732 16580 7744
rect 14507 7704 16580 7732
rect 14507 7701 14519 7704
rect 14461 7695 14519 7701
rect 16574 7692 16580 7704
rect 16632 7692 16638 7744
rect 16684 7732 16712 7828
rect 19886 7760 19892 7812
rect 19944 7800 19950 7812
rect 20073 7803 20131 7809
rect 20073 7800 20085 7803
rect 19944 7772 20085 7800
rect 19944 7760 19950 7772
rect 20073 7769 20085 7772
rect 20119 7800 20131 7803
rect 21560 7800 21588 7831
rect 22830 7828 22836 7840
rect 22888 7828 22894 7880
rect 20119 7772 21588 7800
rect 20119 7769 20131 7772
rect 20073 7763 20131 7769
rect 16853 7735 16911 7741
rect 16853 7732 16865 7735
rect 16684 7704 16865 7732
rect 16853 7701 16865 7704
rect 16899 7701 16911 7735
rect 16853 7695 16911 7701
rect 21358 7692 21364 7744
rect 21416 7732 21422 7744
rect 22281 7735 22339 7741
rect 22281 7732 22293 7735
rect 21416 7704 22293 7732
rect 21416 7692 21422 7704
rect 22281 7701 22293 7704
rect 22327 7701 22339 7735
rect 22281 7695 22339 7701
rect 552 7642 23368 7664
rect 552 7590 3662 7642
rect 3714 7590 3726 7642
rect 3778 7590 3790 7642
rect 3842 7590 3854 7642
rect 3906 7590 3918 7642
rect 3970 7590 23368 7642
rect 552 7568 23368 7590
rect 3142 7488 3148 7540
rect 3200 7528 3206 7540
rect 4617 7531 4675 7537
rect 4617 7528 4629 7531
rect 3200 7500 4629 7528
rect 3200 7488 3206 7500
rect 4617 7497 4629 7500
rect 4663 7497 4675 7531
rect 4617 7491 4675 7497
rect 7374 7488 7380 7540
rect 7432 7488 7438 7540
rect 7926 7488 7932 7540
rect 7984 7488 7990 7540
rect 8386 7488 8392 7540
rect 8444 7488 8450 7540
rect 8573 7531 8631 7537
rect 8573 7497 8585 7531
rect 8619 7497 8631 7531
rect 8573 7491 8631 7497
rect 8202 7420 8208 7472
rect 8260 7460 8266 7472
rect 8588 7460 8616 7491
rect 13262 7488 13268 7540
rect 13320 7488 13326 7540
rect 13998 7488 14004 7540
rect 14056 7488 14062 7540
rect 14274 7488 14280 7540
rect 14332 7488 14338 7540
rect 18782 7488 18788 7540
rect 18840 7488 18846 7540
rect 18969 7531 19027 7537
rect 18969 7497 18981 7531
rect 19015 7528 19027 7531
rect 19245 7531 19303 7537
rect 19245 7528 19257 7531
rect 19015 7500 19257 7528
rect 19015 7497 19027 7500
rect 18969 7491 19027 7497
rect 19245 7497 19257 7500
rect 19291 7497 19303 7531
rect 19245 7491 19303 7497
rect 20714 7488 20720 7540
rect 20772 7488 20778 7540
rect 21358 7488 21364 7540
rect 21416 7488 21422 7540
rect 8260 7432 8616 7460
rect 8260 7420 8266 7432
rect 2866 7352 2872 7404
rect 2924 7392 2930 7404
rect 3234 7392 3240 7404
rect 2924 7364 3240 7392
rect 2924 7352 2930 7364
rect 3234 7352 3240 7364
rect 3292 7352 3298 7404
rect 4706 7352 4712 7404
rect 4764 7352 4770 7404
rect 6914 7352 6920 7404
rect 6972 7392 6978 7404
rect 7009 7395 7067 7401
rect 7009 7392 7021 7395
rect 6972 7364 7021 7392
rect 6972 7352 6978 7364
rect 7009 7361 7021 7364
rect 7055 7361 7067 7395
rect 8220 7392 8248 7420
rect 7009 7355 7067 7361
rect 8128 7364 8248 7392
rect 10781 7395 10839 7401
rect 1673 7327 1731 7333
rect 1673 7293 1685 7327
rect 1719 7324 1731 7327
rect 2884 7324 2912 7352
rect 1719 7296 2912 7324
rect 1719 7293 1731 7296
rect 1673 7287 1731 7293
rect 3050 7284 3056 7336
rect 3108 7284 3114 7336
rect 4724 7324 4752 7352
rect 4890 7324 4896 7336
rect 4724 7296 4896 7324
rect 4890 7284 4896 7296
rect 4948 7284 4954 7336
rect 7101 7327 7159 7333
rect 7101 7293 7113 7327
rect 7147 7324 7159 7327
rect 7190 7324 7196 7336
rect 7147 7296 7196 7324
rect 7147 7293 7159 7296
rect 7101 7287 7159 7293
rect 7190 7284 7196 7296
rect 7248 7284 7254 7336
rect 8128 7333 8156 7364
rect 10781 7361 10793 7395
rect 10827 7392 10839 7395
rect 11606 7392 11612 7404
rect 10827 7364 11612 7392
rect 10827 7361 10839 7364
rect 10781 7355 10839 7361
rect 11606 7352 11612 7364
rect 11664 7352 11670 7404
rect 12802 7352 12808 7404
rect 12860 7352 12866 7404
rect 13630 7352 13636 7404
rect 13688 7352 13694 7404
rect 14458 7352 14464 7404
rect 14516 7352 14522 7404
rect 16850 7392 16856 7404
rect 16040 7364 16856 7392
rect 8113 7327 8171 7333
rect 8113 7293 8125 7327
rect 8159 7293 8171 7327
rect 8113 7287 8171 7293
rect 8202 7284 8208 7336
rect 8260 7284 8266 7336
rect 10686 7284 10692 7336
rect 10744 7284 10750 7336
rect 12897 7327 12955 7333
rect 12897 7293 12909 7327
rect 12943 7324 12955 7327
rect 12986 7324 12992 7336
rect 12943 7296 12992 7324
rect 12943 7293 12955 7296
rect 12897 7287 12955 7293
rect 12986 7284 12992 7296
rect 13044 7284 13050 7336
rect 13725 7327 13783 7333
rect 13725 7293 13737 7327
rect 13771 7324 13783 7327
rect 13814 7324 13820 7336
rect 13771 7296 13820 7324
rect 13771 7293 13783 7296
rect 13725 7287 13783 7293
rect 13814 7284 13820 7296
rect 13872 7284 13878 7336
rect 14550 7284 14556 7336
rect 14608 7284 14614 7336
rect 15562 7284 15568 7336
rect 15620 7324 15626 7336
rect 16040 7333 16068 7364
rect 16850 7352 16856 7364
rect 16908 7352 16914 7404
rect 19426 7392 19432 7404
rect 18340 7364 19432 7392
rect 16025 7327 16083 7333
rect 16025 7324 16037 7327
rect 15620 7296 16037 7324
rect 15620 7284 15626 7296
rect 16025 7293 16037 7296
rect 16071 7293 16083 7327
rect 16025 7287 16083 7293
rect 16209 7327 16267 7333
rect 16209 7293 16221 7327
rect 16255 7324 16267 7327
rect 16482 7324 16488 7336
rect 16255 7296 16488 7324
rect 16255 7293 16267 7296
rect 16209 7287 16267 7293
rect 16482 7284 16488 7296
rect 16540 7284 16546 7336
rect 18340 7333 18368 7364
rect 19426 7352 19432 7364
rect 19484 7392 19490 7404
rect 19886 7392 19892 7404
rect 19484 7364 19656 7392
rect 19484 7352 19490 7364
rect 19628 7333 19656 7364
rect 19720 7364 19892 7392
rect 18325 7327 18383 7333
rect 18325 7293 18337 7327
rect 18371 7293 18383 7327
rect 18325 7287 18383 7293
rect 18509 7327 18567 7333
rect 18509 7293 18521 7327
rect 18555 7324 18567 7327
rect 19613 7327 19671 7333
rect 18555 7296 19472 7324
rect 18555 7293 18567 7296
rect 18509 7287 18567 7293
rect 1940 7259 1998 7265
rect 1940 7225 1952 7259
rect 1986 7256 1998 7259
rect 2130 7256 2136 7268
rect 1986 7228 2136 7256
rect 1986 7225 1998 7228
rect 1940 7219 1998 7225
rect 2130 7216 2136 7228
rect 2188 7216 2194 7268
rect 3068 7256 3096 7284
rect 3482 7259 3540 7265
rect 3482 7256 3494 7259
rect 3068 7228 3494 7256
rect 3482 7225 3494 7228
rect 3528 7225 3540 7259
rect 3482 7219 3540 7225
rect 3694 7216 3700 7268
rect 3752 7256 3758 7268
rect 4709 7259 4767 7265
rect 4709 7256 4721 7259
rect 3752 7228 4721 7256
rect 3752 7216 3758 7228
rect 4709 7225 4721 7228
rect 4755 7225 4767 7259
rect 4709 7219 4767 7225
rect 7650 7216 7656 7268
rect 7708 7256 7714 7268
rect 7929 7259 7987 7265
rect 7929 7256 7941 7259
rect 7708 7228 7941 7256
rect 7708 7216 7714 7228
rect 7929 7225 7941 7228
rect 7975 7256 7987 7259
rect 8757 7259 8815 7265
rect 8757 7256 8769 7259
rect 7975 7228 8769 7256
rect 7975 7225 7987 7228
rect 7929 7219 7987 7225
rect 8757 7225 8769 7228
rect 8803 7225 8815 7259
rect 8757 7219 8815 7225
rect 18417 7259 18475 7265
rect 18417 7225 18429 7259
rect 18463 7256 18475 7259
rect 18937 7259 18995 7265
rect 18937 7256 18949 7259
rect 18463 7228 18949 7256
rect 18463 7225 18475 7228
rect 18417 7219 18475 7225
rect 18937 7225 18949 7228
rect 18983 7225 18995 7259
rect 18937 7219 18995 7225
rect 19150 7216 19156 7268
rect 19208 7216 19214 7268
rect 19444 7265 19472 7296
rect 19613 7293 19625 7327
rect 19659 7293 19671 7327
rect 19613 7287 19671 7293
rect 19429 7259 19487 7265
rect 19429 7225 19441 7259
rect 19475 7256 19487 7259
rect 19720 7256 19748 7364
rect 19886 7352 19892 7364
rect 19944 7352 19950 7404
rect 21910 7392 21916 7404
rect 20824 7364 21916 7392
rect 19794 7284 19800 7336
rect 19852 7324 19858 7336
rect 20073 7327 20131 7333
rect 20073 7324 20085 7327
rect 19852 7296 20085 7324
rect 19852 7284 19858 7296
rect 20073 7293 20085 7296
rect 20119 7293 20131 7327
rect 20073 7287 20131 7293
rect 19475 7228 19748 7256
rect 19889 7259 19947 7265
rect 19475 7225 19487 7228
rect 19429 7219 19487 7225
rect 19889 7225 19901 7259
rect 19935 7256 19947 7259
rect 19978 7256 19984 7268
rect 19935 7228 19984 7256
rect 19935 7225 19947 7228
rect 19889 7219 19947 7225
rect 19978 7216 19984 7228
rect 20036 7216 20042 7268
rect 20701 7259 20759 7265
rect 20701 7225 20713 7259
rect 20747 7256 20759 7259
rect 20824 7256 20852 7364
rect 21910 7352 21916 7364
rect 21968 7352 21974 7404
rect 22186 7352 22192 7404
rect 22244 7392 22250 7404
rect 22370 7392 22376 7404
rect 22244 7364 22376 7392
rect 22244 7352 22250 7364
rect 22370 7352 22376 7364
rect 22428 7352 22434 7404
rect 20990 7284 20996 7336
rect 21048 7284 21054 7336
rect 22462 7284 22468 7336
rect 22520 7284 22526 7336
rect 20747 7228 20852 7256
rect 20901 7259 20959 7265
rect 20747 7225 20759 7228
rect 20701 7219 20759 7225
rect 20901 7225 20913 7259
rect 20947 7256 20959 7259
rect 21818 7256 21824 7268
rect 20947 7228 21824 7256
rect 20947 7225 20959 7228
rect 20901 7219 20959 7225
rect 21818 7216 21824 7228
rect 21876 7216 21882 7268
rect 3053 7191 3111 7197
rect 3053 7157 3065 7191
rect 3099 7188 3111 7191
rect 3326 7188 3332 7200
rect 3099 7160 3332 7188
rect 3099 7157 3111 7160
rect 3053 7151 3111 7157
rect 3326 7148 3332 7160
rect 3384 7188 3390 7200
rect 3602 7188 3608 7200
rect 3384 7160 3608 7188
rect 3384 7148 3390 7160
rect 3602 7148 3608 7160
rect 3660 7148 3666 7200
rect 4798 7148 4804 7200
rect 4856 7188 4862 7200
rect 5077 7191 5135 7197
rect 5077 7188 5089 7191
rect 4856 7160 5089 7188
rect 4856 7148 4862 7160
rect 5077 7157 5089 7160
rect 5123 7157 5135 7191
rect 5077 7151 5135 7157
rect 8202 7148 8208 7200
rect 8260 7188 8266 7200
rect 8547 7191 8605 7197
rect 8547 7188 8559 7191
rect 8260 7160 8559 7188
rect 8260 7148 8266 7160
rect 8547 7157 8559 7160
rect 8593 7157 8605 7191
rect 8547 7151 8605 7157
rect 11057 7191 11115 7197
rect 11057 7157 11069 7191
rect 11103 7188 11115 7191
rect 11606 7188 11612 7200
rect 11103 7160 11612 7188
rect 11103 7157 11115 7160
rect 11057 7151 11115 7157
rect 11606 7148 11612 7160
rect 11664 7148 11670 7200
rect 16206 7148 16212 7200
rect 16264 7148 16270 7200
rect 19334 7148 19340 7200
rect 19392 7188 19398 7200
rect 19705 7191 19763 7197
rect 19705 7188 19717 7191
rect 19392 7160 19717 7188
rect 19392 7148 19398 7160
rect 19705 7157 19717 7160
rect 19751 7157 19763 7191
rect 19705 7151 19763 7157
rect 20530 7148 20536 7200
rect 20588 7148 20594 7200
rect 21266 7148 21272 7200
rect 21324 7188 21330 7200
rect 21361 7191 21419 7197
rect 21361 7188 21373 7191
rect 21324 7160 21373 7188
rect 21324 7148 21330 7160
rect 21361 7157 21373 7160
rect 21407 7157 21419 7191
rect 21361 7151 21419 7157
rect 21542 7148 21548 7200
rect 21600 7148 21606 7200
rect 552 7098 23368 7120
rect 552 7046 4322 7098
rect 4374 7046 4386 7098
rect 4438 7046 4450 7098
rect 4502 7046 4514 7098
rect 4566 7046 4578 7098
rect 4630 7046 23368 7098
rect 552 7024 23368 7046
rect 2130 6944 2136 6996
rect 2188 6944 2194 6996
rect 2301 6987 2359 6993
rect 2301 6953 2313 6987
rect 2347 6984 2359 6987
rect 2406 6984 2412 6996
rect 2347 6956 2412 6984
rect 2347 6953 2359 6956
rect 2301 6947 2359 6953
rect 2406 6944 2412 6956
rect 2464 6944 2470 6996
rect 3050 6944 3056 6996
rect 3108 6984 3114 6996
rect 3145 6987 3203 6993
rect 3145 6984 3157 6987
rect 3108 6956 3157 6984
rect 3108 6944 3114 6956
rect 3145 6953 3157 6956
rect 3191 6953 3203 6987
rect 3145 6947 3203 6953
rect 3237 6987 3295 6993
rect 3237 6953 3249 6987
rect 3283 6984 3295 6987
rect 3694 6984 3700 6996
rect 3283 6956 3700 6984
rect 3283 6953 3295 6956
rect 3237 6947 3295 6953
rect 2501 6919 2559 6925
rect 2501 6885 2513 6919
rect 2547 6916 2559 6919
rect 2774 6916 2780 6928
rect 2547 6888 2780 6916
rect 2547 6885 2559 6888
rect 2501 6879 2559 6885
rect 2774 6876 2780 6888
rect 2832 6916 2838 6928
rect 2961 6919 3019 6925
rect 2961 6916 2973 6919
rect 2832 6888 2973 6916
rect 2832 6876 2838 6888
rect 2961 6885 2973 6888
rect 3007 6885 3019 6919
rect 2961 6879 3019 6885
rect 2593 6851 2651 6857
rect 2593 6817 2605 6851
rect 2639 6848 2651 6851
rect 3252 6848 3280 6947
rect 3694 6944 3700 6956
rect 3752 6944 3758 6996
rect 4249 6987 4307 6993
rect 4249 6953 4261 6987
rect 4295 6984 4307 6987
rect 4890 6984 4896 6996
rect 4295 6956 4896 6984
rect 4295 6953 4307 6956
rect 4249 6947 4307 6953
rect 4890 6944 4896 6956
rect 4948 6944 4954 6996
rect 17497 6987 17555 6993
rect 17497 6953 17509 6987
rect 17543 6953 17555 6987
rect 17497 6947 17555 6953
rect 20993 6987 21051 6993
rect 20993 6953 21005 6987
rect 21039 6984 21051 6987
rect 21450 6984 21456 6996
rect 21039 6956 21456 6984
rect 21039 6953 21051 6956
rect 20993 6947 21051 6953
rect 3418 6925 3424 6928
rect 3405 6919 3424 6925
rect 3405 6885 3417 6919
rect 3405 6879 3424 6885
rect 3418 6876 3424 6879
rect 3476 6876 3482 6928
rect 3602 6876 3608 6928
rect 3660 6876 3666 6928
rect 9766 6876 9772 6928
rect 9824 6916 9830 6928
rect 9824 6888 11284 6916
rect 9824 6876 9830 6888
rect 2639 6820 3280 6848
rect 2639 6817 2651 6820
rect 2593 6811 2651 6817
rect 4798 6808 4804 6860
rect 4856 6848 4862 6860
rect 5362 6851 5420 6857
rect 5362 6848 5374 6851
rect 4856 6820 5374 6848
rect 4856 6808 4862 6820
rect 5362 6817 5374 6820
rect 5408 6817 5420 6851
rect 5362 6811 5420 6817
rect 9585 6851 9643 6857
rect 9585 6817 9597 6851
rect 9631 6848 9643 6851
rect 10042 6848 10048 6860
rect 9631 6820 10048 6848
rect 9631 6817 9643 6820
rect 9585 6811 9643 6817
rect 10042 6808 10048 6820
rect 10100 6808 10106 6860
rect 11146 6808 11152 6860
rect 11204 6808 11210 6860
rect 11256 6848 11284 6888
rect 15562 6876 15568 6928
rect 15620 6876 15626 6928
rect 15749 6919 15807 6925
rect 15749 6885 15761 6919
rect 15795 6916 15807 6919
rect 16482 6916 16488 6928
rect 15795 6888 16488 6916
rect 15795 6885 15807 6888
rect 15749 6879 15807 6885
rect 16482 6876 16488 6888
rect 16540 6916 16546 6928
rect 17512 6916 17540 6947
rect 21450 6944 21456 6956
rect 21508 6944 21514 6996
rect 16540 6888 17540 6916
rect 16540 6876 16546 6888
rect 19978 6876 19984 6928
rect 20036 6916 20042 6928
rect 20809 6919 20867 6925
rect 20809 6916 20821 6919
rect 20036 6888 20821 6916
rect 20036 6876 20042 6888
rect 16390 6857 16396 6860
rect 11609 6851 11667 6857
rect 11609 6848 11621 6851
rect 11256 6820 11621 6848
rect 11609 6817 11621 6820
rect 11655 6817 11667 6851
rect 11609 6811 11667 6817
rect 11885 6851 11943 6857
rect 11885 6817 11897 6851
rect 11931 6817 11943 6851
rect 11885 6811 11943 6817
rect 16384 6811 16396 6857
rect 5626 6740 5632 6792
rect 5684 6740 5690 6792
rect 9490 6740 9496 6792
rect 9548 6740 9554 6792
rect 11054 6740 11060 6792
rect 11112 6740 11118 6792
rect 11701 6783 11759 6789
rect 11701 6780 11713 6783
rect 11164 6752 11713 6780
rect 9953 6715 10011 6721
rect 9953 6681 9965 6715
rect 9999 6712 10011 6715
rect 11164 6712 11192 6752
rect 11701 6749 11713 6752
rect 11747 6749 11759 6783
rect 11701 6743 11759 6749
rect 9999 6684 11192 6712
rect 11517 6715 11575 6721
rect 9999 6681 10011 6684
rect 9953 6675 10011 6681
rect 11517 6681 11529 6715
rect 11563 6712 11575 6715
rect 11900 6712 11928 6811
rect 16390 6808 16396 6811
rect 16448 6808 16454 6860
rect 18322 6808 18328 6860
rect 18380 6808 18386 6860
rect 18598 6857 18604 6860
rect 18592 6811 18604 6857
rect 18598 6808 18604 6811
rect 18656 6808 18662 6860
rect 19886 6808 19892 6860
rect 19944 6808 19950 6860
rect 20088 6857 20116 6888
rect 20809 6885 20821 6888
rect 20855 6885 20867 6919
rect 20809 6879 20867 6885
rect 21542 6876 21548 6928
rect 21600 6916 21606 6928
rect 21698 6919 21756 6925
rect 21698 6916 21710 6919
rect 21600 6888 21710 6916
rect 21600 6876 21606 6888
rect 21698 6885 21710 6888
rect 21744 6885 21756 6919
rect 21698 6879 21756 6885
rect 20073 6851 20131 6857
rect 20073 6817 20085 6851
rect 20119 6817 20131 6851
rect 20073 6811 20131 6817
rect 20165 6851 20223 6857
rect 20165 6817 20177 6851
rect 20211 6848 20223 6851
rect 20254 6848 20260 6860
rect 20211 6820 20260 6848
rect 20211 6817 20223 6820
rect 20165 6811 20223 6817
rect 15930 6740 15936 6792
rect 15988 6780 15994 6792
rect 16117 6783 16175 6789
rect 16117 6780 16129 6783
rect 15988 6752 16129 6780
rect 15988 6740 15994 6752
rect 16117 6749 16129 6752
rect 16163 6749 16175 6783
rect 16117 6743 16175 6749
rect 11563 6684 11928 6712
rect 12069 6715 12127 6721
rect 11563 6681 11575 6684
rect 11517 6675 11575 6681
rect 12069 6681 12081 6715
rect 12115 6712 12127 6715
rect 13906 6712 13912 6724
rect 12115 6684 13912 6712
rect 12115 6681 12127 6684
rect 12069 6675 12127 6681
rect 13906 6672 13912 6684
rect 13964 6672 13970 6724
rect 19702 6672 19708 6724
rect 19760 6712 19766 6724
rect 20088 6712 20116 6811
rect 20254 6808 20260 6820
rect 20312 6848 20318 6860
rect 20625 6851 20683 6857
rect 20625 6848 20637 6851
rect 20312 6820 20637 6848
rect 20312 6808 20318 6820
rect 20625 6817 20637 6820
rect 20671 6817 20683 6851
rect 20625 6811 20683 6817
rect 20717 6851 20775 6857
rect 20717 6817 20729 6851
rect 20763 6817 20775 6851
rect 20717 6811 20775 6817
rect 20732 6780 20760 6811
rect 21174 6808 21180 6860
rect 21232 6848 21238 6860
rect 21453 6851 21511 6857
rect 21453 6848 21465 6851
rect 21232 6820 21465 6848
rect 21232 6808 21238 6820
rect 21453 6817 21465 6820
rect 21499 6817 21511 6851
rect 21453 6811 21511 6817
rect 19760 6684 20116 6712
rect 20180 6752 20760 6780
rect 19760 6672 19766 6684
rect 2314 6604 2320 6656
rect 2372 6604 2378 6656
rect 2958 6604 2964 6656
rect 3016 6604 3022 6656
rect 3234 6604 3240 6656
rect 3292 6644 3298 6656
rect 3421 6647 3479 6653
rect 3421 6644 3433 6647
rect 3292 6616 3433 6644
rect 3292 6604 3298 6616
rect 3421 6613 3433 6616
rect 3467 6613 3479 6647
rect 3421 6607 3479 6613
rect 11606 6604 11612 6656
rect 11664 6604 11670 6656
rect 15933 6647 15991 6653
rect 15933 6613 15945 6647
rect 15979 6644 15991 6647
rect 16114 6644 16120 6656
rect 15979 6616 16120 6644
rect 15979 6613 15991 6616
rect 15933 6607 15991 6613
rect 16114 6604 16120 6616
rect 16172 6604 16178 6656
rect 19978 6604 19984 6656
rect 20036 6644 20042 6656
rect 20180 6653 20208 6752
rect 20898 6740 20904 6792
rect 20956 6780 20962 6792
rect 21266 6780 21272 6792
rect 20956 6752 21272 6780
rect 20956 6740 20962 6752
rect 21266 6740 21272 6752
rect 21324 6740 21330 6792
rect 20441 6715 20499 6721
rect 20441 6681 20453 6715
rect 20487 6712 20499 6715
rect 20714 6712 20720 6724
rect 20487 6684 20720 6712
rect 20487 6681 20499 6684
rect 20441 6675 20499 6681
rect 20714 6672 20720 6684
rect 20772 6672 20778 6724
rect 20165 6647 20223 6653
rect 20165 6644 20177 6647
rect 20036 6616 20177 6644
rect 20036 6604 20042 6616
rect 20165 6613 20177 6616
rect 20211 6613 20223 6647
rect 20165 6607 20223 6613
rect 20349 6647 20407 6653
rect 20349 6613 20361 6647
rect 20395 6644 20407 6647
rect 21266 6644 21272 6656
rect 20395 6616 21272 6644
rect 20395 6613 20407 6616
rect 20349 6607 20407 6613
rect 21266 6604 21272 6616
rect 21324 6604 21330 6656
rect 21818 6604 21824 6656
rect 21876 6644 21882 6656
rect 22833 6647 22891 6653
rect 22833 6644 22845 6647
rect 21876 6616 22845 6644
rect 21876 6604 21882 6616
rect 22833 6613 22845 6616
rect 22879 6613 22891 6647
rect 22833 6607 22891 6613
rect 552 6554 23368 6576
rect 552 6502 3662 6554
rect 3714 6502 3726 6554
rect 3778 6502 3790 6554
rect 3842 6502 3854 6554
rect 3906 6502 3918 6554
rect 3970 6502 23368 6554
rect 552 6480 23368 6502
rect 4617 6443 4675 6449
rect 4617 6409 4629 6443
rect 4663 6440 4675 6443
rect 4706 6440 4712 6452
rect 4663 6412 4712 6440
rect 4663 6409 4675 6412
rect 4617 6403 4675 6409
rect 4706 6400 4712 6412
rect 4764 6400 4770 6452
rect 4798 6400 4804 6452
rect 4856 6400 4862 6452
rect 5721 6443 5779 6449
rect 5721 6409 5733 6443
rect 5767 6440 5779 6443
rect 6089 6443 6147 6449
rect 6089 6440 6101 6443
rect 5767 6412 6101 6440
rect 5767 6409 5779 6412
rect 5721 6403 5779 6409
rect 6089 6409 6101 6412
rect 6135 6409 6147 6443
rect 6089 6403 6147 6409
rect 6457 6443 6515 6449
rect 6457 6409 6469 6443
rect 6503 6440 6515 6443
rect 6917 6443 6975 6449
rect 6917 6440 6929 6443
rect 6503 6412 6929 6440
rect 6503 6409 6515 6412
rect 6457 6403 6515 6409
rect 6917 6409 6929 6412
rect 6963 6409 6975 6443
rect 6917 6403 6975 6409
rect 13814 6400 13820 6452
rect 13872 6440 13878 6452
rect 14274 6440 14280 6452
rect 13872 6412 14280 6440
rect 13872 6400 13878 6412
rect 14274 6400 14280 6412
rect 14332 6400 14338 6452
rect 14645 6443 14703 6449
rect 14645 6409 14657 6443
rect 14691 6440 14703 6443
rect 15562 6440 15568 6452
rect 14691 6412 15568 6440
rect 14691 6409 14703 6412
rect 14645 6403 14703 6409
rect 15562 6400 15568 6412
rect 15620 6400 15626 6452
rect 16206 6400 16212 6452
rect 16264 6400 16270 6452
rect 16390 6400 16396 6452
rect 16448 6400 16454 6452
rect 18598 6400 18604 6452
rect 18656 6440 18662 6452
rect 18693 6443 18751 6449
rect 18693 6440 18705 6443
rect 18656 6412 18705 6440
rect 18656 6400 18662 6412
rect 18693 6409 18705 6412
rect 18739 6409 18751 6443
rect 18693 6403 18751 6409
rect 18877 6443 18935 6449
rect 18877 6409 18889 6443
rect 18923 6440 18935 6443
rect 19150 6440 19156 6452
rect 18923 6412 19156 6440
rect 18923 6409 18935 6412
rect 18877 6403 18935 6409
rect 19150 6400 19156 6412
rect 19208 6400 19214 6452
rect 19337 6443 19395 6449
rect 19337 6409 19349 6443
rect 19383 6440 19395 6443
rect 19426 6440 19432 6452
rect 19383 6412 19432 6440
rect 19383 6409 19395 6412
rect 19337 6403 19395 6409
rect 19426 6400 19432 6412
rect 19484 6400 19490 6452
rect 19794 6400 19800 6452
rect 19852 6400 19858 6452
rect 19978 6400 19984 6452
rect 20036 6400 20042 6452
rect 20898 6400 20904 6452
rect 20956 6440 20962 6452
rect 21138 6443 21196 6449
rect 21138 6440 21150 6443
rect 20956 6412 21150 6440
rect 20956 6400 20962 6412
rect 21138 6409 21150 6412
rect 21184 6409 21196 6443
rect 22094 6440 22100 6452
rect 21138 6403 21196 6409
rect 21284 6412 22100 6440
rect 4246 6332 4252 6384
rect 4304 6332 4310 6384
rect 5810 6332 5816 6384
rect 5868 6372 5874 6384
rect 6822 6372 6828 6384
rect 5868 6344 6828 6372
rect 5868 6332 5874 6344
rect 6822 6332 6828 6344
rect 6880 6372 6886 6384
rect 6880 6344 7328 6372
rect 6880 6332 6886 6344
rect 6730 6304 6736 6316
rect 6288 6276 6736 6304
rect 5810 6196 5816 6248
rect 5868 6236 5874 6248
rect 5997 6239 6055 6245
rect 5997 6236 6009 6239
rect 5868 6208 6009 6236
rect 5868 6196 5874 6208
rect 5997 6205 6009 6208
rect 6043 6205 6055 6239
rect 5997 6199 6055 6205
rect 6181 6239 6239 6245
rect 6181 6205 6193 6239
rect 6227 6230 6239 6239
rect 6288 6230 6316 6276
rect 6730 6264 6736 6276
rect 6788 6264 6794 6316
rect 6227 6205 6316 6230
rect 6181 6202 6316 6205
rect 6181 6199 6239 6202
rect 6546 6196 6552 6248
rect 6604 6236 6610 6248
rect 6825 6239 6883 6245
rect 6825 6236 6837 6239
rect 6604 6208 6837 6236
rect 6604 6196 6610 6208
rect 6825 6205 6837 6208
rect 6871 6205 6883 6239
rect 6825 6199 6883 6205
rect 7101 6239 7159 6245
rect 7101 6205 7113 6239
rect 7147 6236 7159 6239
rect 7190 6236 7196 6248
rect 7147 6208 7196 6236
rect 7147 6205 7159 6208
rect 7101 6199 7159 6205
rect 5905 6171 5963 6177
rect 5905 6168 5917 6171
rect 4632 6140 5917 6168
rect 3510 6060 3516 6112
rect 3568 6100 3574 6112
rect 4632 6109 4660 6140
rect 5905 6137 5917 6140
rect 5951 6168 5963 6171
rect 6840 6168 6868 6199
rect 7190 6196 7196 6208
rect 7248 6196 7254 6248
rect 7300 6245 7328 6344
rect 11974 6332 11980 6384
rect 12032 6372 12038 6384
rect 21284 6372 21312 6412
rect 22094 6400 22100 6412
rect 22152 6400 22158 6452
rect 12032 6344 21312 6372
rect 12032 6332 12038 6344
rect 19245 6307 19303 6313
rect 19245 6273 19257 6307
rect 19291 6304 19303 6307
rect 19426 6304 19432 6316
rect 19291 6276 19432 6304
rect 19291 6273 19303 6276
rect 19245 6267 19303 6273
rect 19426 6264 19432 6276
rect 19484 6264 19490 6316
rect 19702 6264 19708 6316
rect 19760 6264 19766 6316
rect 20530 6264 20536 6316
rect 20588 6304 20594 6316
rect 20809 6307 20867 6313
rect 20809 6304 20821 6307
rect 20588 6276 20821 6304
rect 20588 6264 20594 6276
rect 20809 6273 20821 6276
rect 20855 6273 20867 6307
rect 20809 6267 20867 6273
rect 21192 6276 21588 6304
rect 7285 6239 7343 6245
rect 7285 6205 7297 6239
rect 7331 6205 7343 6239
rect 7285 6199 7343 6205
rect 7374 6196 7380 6248
rect 7432 6196 7438 6248
rect 7650 6196 7656 6248
rect 7708 6196 7714 6248
rect 14369 6239 14427 6245
rect 14369 6205 14381 6239
rect 14415 6236 14427 6239
rect 14550 6236 14556 6248
rect 14415 6208 14556 6236
rect 14415 6205 14427 6208
rect 14369 6199 14427 6205
rect 14550 6196 14556 6208
rect 14608 6236 14614 6248
rect 14608 6208 14964 6236
rect 14608 6196 14614 6208
rect 14936 6180 14964 6208
rect 19334 6196 19340 6248
rect 19392 6196 19398 6248
rect 19521 6239 19579 6245
rect 19521 6205 19533 6239
rect 19567 6236 19579 6239
rect 19794 6236 19800 6248
rect 19567 6208 19800 6236
rect 19567 6205 19579 6208
rect 19521 6199 19579 6205
rect 19794 6196 19800 6208
rect 19852 6196 19858 6248
rect 20548 6236 20576 6264
rect 20088 6208 20576 6236
rect 20717 6239 20775 6245
rect 7469 6171 7527 6177
rect 7469 6168 7481 6171
rect 5951 6140 6500 6168
rect 6840 6140 7481 6168
rect 5951 6137 5963 6140
rect 5905 6131 5963 6137
rect 6472 6112 6500 6140
rect 7469 6137 7481 6140
rect 7515 6137 7527 6171
rect 7469 6131 7527 6137
rect 12986 6128 12992 6180
rect 13044 6168 13050 6180
rect 13633 6171 13691 6177
rect 13633 6168 13645 6171
rect 13044 6140 13645 6168
rect 13044 6128 13050 6140
rect 13633 6137 13645 6140
rect 13679 6168 13691 6171
rect 13722 6168 13728 6180
rect 13679 6140 13728 6168
rect 13679 6137 13691 6140
rect 13633 6131 13691 6137
rect 13722 6128 13728 6140
rect 13780 6168 13786 6180
rect 14093 6171 14151 6177
rect 14093 6168 14105 6171
rect 13780 6140 14105 6168
rect 13780 6128 13786 6140
rect 14093 6137 14105 6140
rect 14139 6137 14151 6171
rect 14737 6171 14795 6177
rect 14737 6168 14749 6171
rect 14093 6131 14151 6137
rect 14200 6140 14749 6168
rect 4617 6103 4675 6109
rect 4617 6100 4629 6103
rect 3568 6072 4629 6100
rect 3568 6060 3574 6072
rect 4617 6069 4629 6072
rect 4663 6069 4675 6103
rect 4617 6063 4675 6069
rect 5534 6060 5540 6112
rect 5592 6060 5598 6112
rect 5718 6109 5724 6112
rect 5705 6103 5724 6109
rect 5705 6069 5717 6103
rect 5705 6063 5724 6069
rect 5718 6060 5724 6063
rect 5776 6060 5782 6112
rect 6273 6103 6331 6109
rect 6273 6069 6285 6103
rect 6319 6100 6331 6103
rect 6362 6100 6368 6112
rect 6319 6072 6368 6100
rect 6319 6069 6331 6072
rect 6273 6063 6331 6069
rect 6362 6060 6368 6072
rect 6420 6060 6426 6112
rect 6454 6060 6460 6112
rect 6512 6060 6518 6112
rect 6730 6060 6736 6112
rect 6788 6100 6794 6112
rect 7374 6100 7380 6112
rect 6788 6072 7380 6100
rect 6788 6060 6794 6072
rect 7374 6060 7380 6072
rect 7432 6060 7438 6112
rect 7837 6103 7895 6109
rect 7837 6069 7849 6103
rect 7883 6100 7895 6103
rect 8018 6100 8024 6112
rect 7883 6072 8024 6100
rect 7883 6069 7895 6072
rect 7837 6063 7895 6069
rect 8018 6060 8024 6072
rect 8076 6060 8082 6112
rect 13354 6060 13360 6112
rect 13412 6100 13418 6112
rect 13833 6103 13891 6109
rect 13833 6100 13845 6103
rect 13412 6072 13845 6100
rect 13412 6060 13418 6072
rect 13833 6069 13845 6072
rect 13879 6069 13891 6103
rect 13833 6063 13891 6069
rect 13998 6060 14004 6112
rect 14056 6100 14062 6112
rect 14200 6100 14228 6140
rect 14737 6137 14749 6140
rect 14783 6137 14795 6171
rect 14737 6131 14795 6137
rect 14918 6128 14924 6180
rect 14976 6128 14982 6180
rect 16022 6128 16028 6180
rect 16080 6128 16086 6180
rect 16114 6128 16120 6180
rect 16172 6168 16178 6180
rect 16225 6171 16283 6177
rect 16225 6168 16237 6171
rect 16172 6140 16237 6168
rect 16172 6128 16178 6140
rect 16225 6137 16237 6140
rect 16271 6137 16283 6171
rect 16225 6131 16283 6137
rect 18877 6171 18935 6177
rect 18877 6137 18889 6171
rect 18923 6168 18935 6171
rect 19352 6168 19380 6196
rect 18923 6140 19380 6168
rect 19965 6171 20023 6177
rect 18923 6137 18935 6140
rect 18877 6131 18935 6137
rect 19965 6137 19977 6171
rect 20011 6168 20023 6171
rect 20088 6168 20116 6208
rect 20717 6205 20729 6239
rect 20763 6236 20775 6239
rect 21082 6236 21088 6248
rect 20763 6208 21088 6236
rect 20763 6205 20775 6208
rect 20717 6199 20775 6205
rect 21082 6196 21088 6208
rect 21140 6196 21146 6248
rect 20011 6140 20116 6168
rect 20165 6171 20223 6177
rect 20011 6137 20023 6140
rect 19965 6131 20023 6137
rect 20165 6137 20177 6171
rect 20211 6168 20223 6171
rect 20254 6168 20260 6180
rect 20211 6140 20260 6168
rect 20211 6137 20223 6140
rect 20165 6131 20223 6137
rect 20254 6128 20260 6140
rect 20312 6128 20318 6180
rect 20533 6171 20591 6177
rect 20533 6137 20545 6171
rect 20579 6168 20591 6171
rect 20806 6168 20812 6180
rect 20579 6140 20812 6168
rect 20579 6137 20591 6140
rect 20533 6131 20591 6137
rect 14056 6072 14228 6100
rect 14056 6060 14062 6072
rect 14274 6060 14280 6112
rect 14332 6060 14338 6112
rect 14461 6103 14519 6109
rect 14461 6069 14473 6103
rect 14507 6100 14519 6103
rect 14550 6100 14556 6112
rect 14507 6072 14556 6100
rect 14507 6069 14519 6072
rect 14461 6063 14519 6069
rect 14550 6060 14556 6072
rect 14608 6060 14614 6112
rect 15105 6103 15163 6109
rect 15105 6069 15117 6103
rect 15151 6100 15163 6103
rect 15194 6100 15200 6112
rect 15151 6072 15200 6100
rect 15151 6069 15163 6072
rect 15105 6063 15163 6069
rect 15194 6060 15200 6072
rect 15252 6060 15258 6112
rect 15930 6060 15936 6112
rect 15988 6100 15994 6112
rect 16482 6100 16488 6112
rect 15988 6072 16488 6100
rect 15988 6060 15994 6072
rect 16482 6060 16488 6072
rect 16540 6100 16546 6112
rect 20548 6100 20576 6131
rect 20806 6128 20812 6140
rect 20864 6128 20870 6180
rect 16540 6072 20576 6100
rect 21100 6100 21128 6196
rect 21192 6177 21220 6276
rect 21453 6239 21511 6245
rect 21453 6236 21465 6239
rect 21284 6208 21465 6236
rect 21177 6171 21235 6177
rect 21177 6137 21189 6171
rect 21223 6137 21235 6171
rect 21177 6131 21235 6137
rect 21284 6100 21312 6208
rect 21453 6205 21465 6208
rect 21499 6205 21511 6239
rect 21560 6236 21588 6276
rect 22554 6236 22560 6248
rect 21560 6208 22560 6236
rect 21453 6199 21511 6205
rect 22554 6196 22560 6208
rect 22612 6196 22618 6248
rect 21698 6171 21756 6177
rect 21698 6168 21710 6171
rect 21376 6140 21710 6168
rect 21376 6109 21404 6140
rect 21698 6137 21710 6140
rect 21744 6137 21756 6171
rect 21698 6131 21756 6137
rect 21100 6072 21312 6100
rect 21361 6103 21419 6109
rect 16540 6060 16546 6072
rect 21361 6069 21373 6103
rect 21407 6069 21419 6103
rect 21361 6063 21419 6069
rect 22830 6060 22836 6112
rect 22888 6060 22894 6112
rect 552 6010 23368 6032
rect 552 5958 4322 6010
rect 4374 5958 4386 6010
rect 4438 5958 4450 6010
rect 4502 5958 4514 6010
rect 4566 5958 4578 6010
rect 4630 5958 23368 6010
rect 552 5936 23368 5958
rect 5629 5899 5687 5905
rect 5629 5865 5641 5899
rect 5675 5896 5687 5899
rect 5718 5896 5724 5908
rect 5675 5868 5724 5896
rect 5675 5865 5687 5868
rect 5629 5859 5687 5865
rect 5718 5856 5724 5868
rect 5776 5856 5782 5908
rect 7190 5856 7196 5908
rect 7248 5896 7254 5908
rect 7469 5899 7527 5905
rect 7469 5896 7481 5899
rect 7248 5868 7481 5896
rect 7248 5856 7254 5868
rect 7469 5865 7481 5868
rect 7515 5865 7527 5899
rect 7469 5859 7527 5865
rect 7561 5899 7619 5905
rect 7561 5865 7573 5899
rect 7607 5896 7619 5899
rect 7650 5896 7656 5908
rect 7607 5868 7656 5896
rect 7607 5865 7619 5868
rect 7561 5859 7619 5865
rect 7650 5856 7656 5868
rect 7708 5856 7714 5908
rect 9398 5896 9404 5908
rect 9140 5868 9404 5896
rect 4246 5788 4252 5840
rect 4304 5828 4310 5840
rect 5261 5831 5319 5837
rect 5261 5828 5273 5831
rect 4304 5800 5273 5828
rect 4304 5788 4310 5800
rect 5261 5797 5273 5800
rect 5307 5797 5319 5831
rect 5261 5791 5319 5797
rect 5445 5831 5503 5837
rect 5445 5797 5457 5831
rect 5491 5828 5503 5831
rect 5810 5828 5816 5840
rect 5491 5800 5816 5828
rect 5491 5797 5503 5800
rect 5445 5791 5503 5797
rect 5276 5760 5304 5791
rect 5810 5788 5816 5800
rect 5868 5788 5874 5840
rect 6730 5828 6736 5840
rect 6196 5800 6736 5828
rect 6196 5760 6224 5800
rect 6730 5788 6736 5800
rect 6788 5788 6794 5840
rect 6362 5769 6368 5772
rect 6356 5760 6368 5769
rect 5276 5732 6224 5760
rect 6323 5732 6368 5760
rect 6356 5723 6368 5732
rect 6362 5720 6368 5723
rect 6420 5720 6426 5772
rect 8294 5720 8300 5772
rect 8352 5760 8358 5772
rect 8674 5763 8732 5769
rect 8674 5760 8686 5763
rect 8352 5732 8686 5760
rect 8352 5720 8358 5732
rect 8674 5729 8686 5732
rect 8720 5729 8732 5763
rect 8674 5723 8732 5729
rect 8846 5720 8852 5772
rect 8904 5760 8910 5772
rect 9140 5769 9168 5868
rect 9398 5856 9404 5868
rect 9456 5896 9462 5908
rect 9456 5868 11100 5896
rect 9456 5856 9462 5868
rect 10042 5828 10048 5840
rect 9324 5800 10048 5828
rect 9324 5769 9352 5800
rect 10042 5788 10048 5800
rect 10100 5788 10106 5840
rect 8941 5763 8999 5769
rect 8941 5760 8953 5763
rect 8904 5732 8953 5760
rect 8904 5720 8910 5732
rect 8941 5729 8953 5732
rect 8987 5729 8999 5763
rect 8941 5723 8999 5729
rect 9125 5763 9183 5769
rect 9125 5729 9137 5763
rect 9171 5729 9183 5763
rect 9125 5723 9183 5729
rect 9309 5763 9367 5769
rect 9309 5729 9321 5763
rect 9355 5729 9367 5763
rect 9309 5723 9367 5729
rect 5626 5652 5632 5704
rect 5684 5692 5690 5704
rect 6089 5695 6147 5701
rect 6089 5692 6101 5695
rect 5684 5664 6101 5692
rect 5684 5652 5690 5664
rect 6089 5661 6101 5664
rect 6135 5661 6147 5695
rect 6089 5655 6147 5661
rect 8956 5624 8984 5723
rect 9858 5720 9864 5772
rect 9916 5720 9922 5772
rect 10152 5769 10180 5868
rect 10226 5788 10232 5840
rect 10284 5828 10290 5840
rect 10965 5831 11023 5837
rect 10965 5828 10977 5831
rect 10284 5800 10977 5828
rect 10284 5788 10290 5800
rect 10965 5797 10977 5800
rect 11011 5797 11023 5831
rect 11072 5828 11100 5868
rect 11146 5856 11152 5908
rect 11204 5896 11210 5908
rect 11241 5899 11299 5905
rect 11241 5896 11253 5899
rect 11204 5868 11253 5896
rect 11204 5856 11210 5868
rect 11241 5865 11253 5868
rect 11287 5865 11299 5899
rect 11241 5859 11299 5865
rect 11974 5856 11980 5908
rect 12032 5856 12038 5908
rect 13722 5856 13728 5908
rect 13780 5896 13786 5908
rect 14461 5899 14519 5905
rect 14461 5896 14473 5899
rect 13780 5868 14473 5896
rect 13780 5856 13786 5868
rect 14461 5865 14473 5868
rect 14507 5865 14519 5899
rect 14461 5859 14519 5865
rect 19978 5856 19984 5908
rect 20036 5856 20042 5908
rect 20254 5856 20260 5908
rect 20312 5896 20318 5908
rect 20441 5899 20499 5905
rect 20441 5896 20453 5899
rect 20312 5868 20453 5896
rect 20312 5856 20318 5868
rect 20441 5865 20453 5868
rect 20487 5865 20499 5899
rect 20441 5859 20499 5865
rect 20990 5856 20996 5908
rect 21048 5896 21054 5908
rect 21729 5899 21787 5905
rect 21729 5896 21741 5899
rect 21048 5868 21741 5896
rect 21048 5856 21054 5868
rect 21729 5865 21741 5868
rect 21775 5896 21787 5899
rect 21775 5868 22232 5896
rect 21775 5865 21787 5868
rect 21729 5859 21787 5865
rect 11333 5831 11391 5837
rect 11333 5828 11345 5831
rect 11072 5800 11345 5828
rect 10965 5791 11023 5797
rect 11333 5797 11345 5800
rect 11379 5797 11391 5831
rect 11333 5791 11391 5797
rect 12526 5788 12532 5840
rect 12584 5828 12590 5840
rect 13633 5831 13691 5837
rect 13633 5828 13645 5831
rect 12584 5800 13645 5828
rect 12584 5788 12590 5800
rect 13633 5797 13645 5800
rect 13679 5828 13691 5831
rect 15197 5831 15255 5837
rect 15197 5828 15209 5831
rect 13679 5800 15209 5828
rect 13679 5797 13691 5800
rect 13633 5791 13691 5797
rect 15197 5797 15209 5800
rect 15243 5828 15255 5831
rect 15378 5828 15384 5840
rect 15243 5800 15384 5828
rect 15243 5797 15255 5800
rect 15197 5791 15255 5797
rect 15378 5788 15384 5800
rect 15436 5828 15442 5840
rect 16022 5828 16028 5840
rect 15436 5800 16028 5828
rect 15436 5788 15442 5800
rect 16022 5788 16028 5800
rect 16080 5788 16086 5840
rect 19702 5828 19708 5840
rect 18616 5800 19708 5828
rect 10137 5763 10195 5769
rect 10137 5729 10149 5763
rect 10183 5729 10195 5763
rect 10137 5723 10195 5729
rect 10413 5763 10471 5769
rect 10413 5729 10425 5763
rect 10459 5760 10471 5763
rect 10686 5760 10692 5772
rect 10459 5732 10692 5760
rect 10459 5729 10471 5732
rect 10413 5723 10471 5729
rect 10686 5720 10692 5732
rect 10744 5760 10750 5772
rect 11149 5763 11207 5769
rect 11149 5760 11161 5763
rect 10744 5732 11161 5760
rect 10744 5720 10750 5732
rect 11149 5729 11161 5732
rect 11195 5729 11207 5763
rect 11149 5723 11207 5729
rect 12986 5720 12992 5772
rect 13044 5720 13050 5772
rect 13173 5763 13231 5769
rect 13173 5729 13185 5763
rect 13219 5729 13231 5763
rect 13173 5723 13231 5729
rect 9876 5692 9904 5720
rect 11422 5692 11428 5704
rect 9876 5664 11428 5692
rect 11422 5652 11428 5664
rect 11480 5652 11486 5704
rect 11517 5695 11575 5701
rect 11517 5661 11529 5695
rect 11563 5692 11575 5695
rect 11609 5695 11667 5701
rect 11609 5692 11621 5695
rect 11563 5664 11621 5692
rect 11563 5661 11575 5664
rect 11517 5655 11575 5661
rect 11609 5661 11621 5664
rect 11655 5692 11667 5695
rect 13188 5692 13216 5723
rect 13998 5720 14004 5772
rect 14056 5720 14062 5772
rect 14274 5720 14280 5772
rect 14332 5720 14338 5772
rect 14550 5720 14556 5772
rect 14608 5720 14614 5772
rect 14829 5763 14887 5769
rect 14829 5729 14841 5763
rect 14875 5760 14887 5763
rect 15562 5760 15568 5772
rect 14875 5732 15568 5760
rect 14875 5729 14887 5732
rect 14829 5723 14887 5729
rect 15562 5720 15568 5732
rect 15620 5720 15626 5772
rect 18322 5720 18328 5772
rect 18380 5760 18386 5772
rect 18616 5769 18644 5800
rect 19702 5788 19708 5800
rect 19760 5788 19766 5840
rect 18874 5769 18880 5772
rect 18601 5763 18659 5769
rect 18601 5760 18613 5763
rect 18380 5732 18613 5760
rect 18380 5720 18386 5732
rect 18601 5729 18613 5732
rect 18647 5729 18659 5763
rect 18601 5723 18659 5729
rect 18868 5723 18880 5769
rect 18874 5720 18880 5723
rect 18932 5720 18938 5772
rect 19996 5760 20024 5856
rect 22204 5837 22232 5868
rect 22554 5856 22560 5908
rect 22612 5856 22618 5908
rect 22189 5831 22247 5837
rect 21836 5800 22048 5828
rect 21836 5772 21864 5800
rect 20257 5763 20315 5769
rect 20257 5760 20269 5763
rect 19996 5732 20269 5760
rect 20257 5729 20269 5732
rect 20303 5729 20315 5763
rect 20257 5723 20315 5729
rect 20346 5720 20352 5772
rect 20404 5760 20410 5772
rect 20533 5763 20591 5769
rect 20533 5760 20545 5763
rect 20404 5732 20545 5760
rect 20404 5720 20410 5732
rect 20533 5729 20545 5732
rect 20579 5760 20591 5763
rect 20622 5760 20628 5772
rect 20579 5732 20628 5760
rect 20579 5729 20591 5732
rect 20533 5723 20591 5729
rect 20622 5720 20628 5732
rect 20680 5720 20686 5772
rect 21266 5720 21272 5772
rect 21324 5720 21330 5772
rect 21453 5763 21511 5769
rect 21453 5729 21465 5763
rect 21499 5760 21511 5763
rect 21818 5760 21824 5772
rect 21499 5732 21824 5760
rect 21499 5729 21511 5732
rect 21453 5723 21511 5729
rect 21818 5720 21824 5732
rect 21876 5720 21882 5772
rect 21910 5720 21916 5772
rect 21968 5720 21974 5772
rect 22020 5769 22048 5800
rect 22189 5797 22201 5831
rect 22235 5797 22247 5831
rect 22189 5791 22247 5797
rect 22005 5763 22063 5769
rect 22005 5729 22017 5763
rect 22051 5729 22063 5763
rect 22005 5723 22063 5729
rect 22373 5763 22431 5769
rect 22373 5729 22385 5763
rect 22419 5760 22431 5763
rect 22830 5760 22836 5772
rect 22419 5732 22836 5760
rect 22419 5729 22431 5732
rect 22373 5723 22431 5729
rect 13354 5692 13360 5704
rect 11655 5664 13360 5692
rect 11655 5661 11667 5664
rect 11609 5655 11667 5661
rect 13354 5652 13360 5664
rect 13412 5692 13418 5704
rect 14568 5692 14596 5720
rect 13412 5664 14596 5692
rect 13412 5652 13418 5664
rect 20714 5652 20720 5704
rect 20772 5692 20778 5704
rect 22388 5692 22416 5723
rect 22830 5720 22836 5732
rect 22888 5720 22894 5772
rect 20772 5664 22416 5692
rect 20772 5652 20778 5664
rect 10045 5627 10103 5633
rect 10045 5624 10057 5627
rect 8956 5596 10057 5624
rect 10045 5593 10057 5596
rect 10091 5593 10103 5627
rect 10045 5587 10103 5593
rect 13449 5627 13507 5633
rect 13449 5593 13461 5627
rect 13495 5624 13507 5627
rect 13814 5624 13820 5636
rect 13495 5596 13820 5624
rect 13495 5593 13507 5596
rect 13449 5587 13507 5593
rect 13814 5584 13820 5596
rect 13872 5584 13878 5636
rect 8754 5516 8760 5568
rect 8812 5556 8818 5568
rect 9217 5559 9275 5565
rect 9217 5556 9229 5559
rect 8812 5528 9229 5556
rect 8812 5516 8818 5528
rect 9217 5525 9229 5528
rect 9263 5525 9275 5559
rect 9217 5519 9275 5525
rect 10318 5516 10324 5568
rect 10376 5556 10382 5568
rect 10597 5559 10655 5565
rect 10597 5556 10609 5559
rect 10376 5528 10609 5556
rect 10376 5516 10382 5528
rect 10597 5525 10609 5528
rect 10643 5525 10655 5559
rect 10597 5519 10655 5525
rect 11974 5516 11980 5568
rect 12032 5516 12038 5568
rect 12066 5516 12072 5568
rect 12124 5556 12130 5568
rect 12161 5559 12219 5565
rect 12161 5556 12173 5559
rect 12124 5528 12173 5556
rect 12124 5516 12130 5528
rect 12161 5525 12173 5528
rect 12207 5525 12219 5559
rect 12161 5519 12219 5525
rect 12710 5516 12716 5568
rect 12768 5556 12774 5568
rect 13081 5559 13139 5565
rect 13081 5556 13093 5559
rect 12768 5528 13093 5556
rect 12768 5516 12774 5528
rect 13081 5525 13093 5528
rect 13127 5525 13139 5559
rect 13081 5519 13139 5525
rect 13633 5559 13691 5565
rect 13633 5525 13645 5559
rect 13679 5556 13691 5559
rect 14093 5559 14151 5565
rect 14093 5556 14105 5559
rect 13679 5528 14105 5556
rect 13679 5525 13691 5528
rect 13633 5519 13691 5525
rect 14093 5525 14105 5528
rect 14139 5525 14151 5559
rect 14093 5519 14151 5525
rect 15194 5516 15200 5568
rect 15252 5516 15258 5568
rect 15378 5516 15384 5568
rect 15436 5516 15442 5568
rect 20070 5516 20076 5568
rect 20128 5516 20134 5568
rect 21453 5559 21511 5565
rect 21453 5525 21465 5559
rect 21499 5556 21511 5559
rect 21560 5556 21588 5664
rect 21637 5627 21695 5633
rect 21637 5593 21649 5627
rect 21683 5624 21695 5627
rect 22278 5624 22284 5636
rect 21683 5596 22284 5624
rect 21683 5593 21695 5596
rect 21637 5587 21695 5593
rect 22278 5584 22284 5596
rect 22336 5584 22342 5636
rect 21499 5528 21588 5556
rect 21499 5525 21511 5528
rect 21453 5519 21511 5525
rect 552 5466 23368 5488
rect 552 5414 3662 5466
rect 3714 5414 3726 5466
rect 3778 5414 3790 5466
rect 3842 5414 3854 5466
rect 3906 5414 3918 5466
rect 3970 5414 23368 5466
rect 552 5392 23368 5414
rect 2685 5355 2743 5361
rect 2685 5321 2697 5355
rect 2731 5352 2743 5355
rect 2774 5352 2780 5364
rect 2731 5324 2780 5352
rect 2731 5321 2743 5324
rect 2685 5315 2743 5321
rect 2774 5312 2780 5324
rect 2832 5352 2838 5364
rect 3510 5352 3516 5364
rect 2832 5324 3516 5352
rect 2832 5312 2838 5324
rect 3510 5312 3516 5324
rect 3568 5312 3574 5364
rect 5626 5352 5632 5364
rect 5460 5324 5632 5352
rect 3053 5287 3111 5293
rect 3053 5253 3065 5287
rect 3099 5284 3111 5287
rect 3418 5284 3424 5296
rect 3099 5256 3424 5284
rect 3099 5253 3111 5256
rect 3053 5247 3111 5253
rect 3418 5244 3424 5256
rect 3476 5284 3482 5296
rect 3878 5284 3884 5296
rect 3476 5256 3884 5284
rect 3476 5244 3482 5256
rect 3878 5244 3884 5256
rect 3936 5244 3942 5296
rect 2866 5108 2872 5160
rect 2924 5148 2930 5160
rect 5460 5157 5488 5324
rect 5626 5312 5632 5324
rect 5684 5312 5690 5364
rect 6822 5312 6828 5364
rect 6880 5352 6886 5364
rect 6880 5312 6914 5352
rect 8018 5312 8024 5364
rect 8076 5312 8082 5364
rect 8205 5355 8263 5361
rect 8205 5321 8217 5355
rect 8251 5352 8263 5355
rect 8294 5352 8300 5364
rect 8251 5324 8300 5352
rect 8251 5321 8263 5324
rect 8205 5315 8263 5321
rect 8294 5312 8300 5324
rect 8352 5312 8358 5364
rect 8754 5312 8760 5364
rect 8812 5312 8818 5364
rect 10686 5312 10692 5364
rect 10744 5352 10750 5364
rect 10873 5355 10931 5361
rect 10873 5352 10885 5355
rect 10744 5324 10885 5352
rect 10744 5312 10750 5324
rect 10873 5321 10885 5324
rect 10919 5321 10931 5355
rect 10873 5315 10931 5321
rect 10965 5355 11023 5361
rect 10965 5321 10977 5355
rect 11011 5352 11023 5355
rect 11146 5352 11152 5364
rect 11011 5324 11152 5352
rect 11011 5321 11023 5324
rect 10965 5315 11023 5321
rect 11146 5312 11152 5324
rect 11204 5312 11210 5364
rect 12710 5312 12716 5364
rect 12768 5312 12774 5364
rect 14918 5312 14924 5364
rect 14976 5352 14982 5364
rect 15105 5355 15163 5361
rect 15105 5352 15117 5355
rect 14976 5324 15117 5352
rect 14976 5312 14982 5324
rect 15105 5321 15117 5324
rect 15151 5321 15163 5355
rect 15105 5315 15163 5321
rect 18785 5355 18843 5361
rect 18785 5321 18797 5355
rect 18831 5352 18843 5355
rect 18874 5352 18880 5364
rect 18831 5324 18880 5352
rect 18831 5321 18843 5324
rect 18785 5315 18843 5321
rect 18874 5312 18880 5324
rect 18932 5312 18938 5364
rect 18969 5355 19027 5361
rect 18969 5321 18981 5355
rect 19015 5352 19027 5355
rect 19150 5352 19156 5364
rect 19015 5324 19156 5352
rect 19015 5321 19027 5324
rect 18969 5315 19027 5321
rect 19150 5312 19156 5324
rect 19208 5312 19214 5364
rect 20806 5312 20812 5364
rect 20864 5352 20870 5364
rect 21729 5355 21787 5361
rect 21729 5352 21741 5355
rect 20864 5324 21741 5352
rect 20864 5312 20870 5324
rect 21729 5321 21741 5324
rect 21775 5321 21787 5355
rect 21729 5315 21787 5321
rect 6886 5284 6914 5312
rect 7009 5287 7067 5293
rect 7009 5284 7021 5287
rect 6886 5256 7021 5284
rect 7009 5253 7021 5256
rect 7055 5253 7067 5287
rect 7009 5247 7067 5253
rect 7561 5287 7619 5293
rect 7561 5253 7573 5287
rect 7607 5284 7619 5287
rect 7607 5256 7696 5284
rect 7607 5253 7619 5256
rect 7561 5247 7619 5253
rect 5445 5151 5503 5157
rect 5445 5148 5457 5151
rect 2924 5120 5457 5148
rect 2924 5108 2930 5120
rect 5445 5117 5457 5120
rect 5491 5117 5503 5151
rect 5445 5111 5503 5117
rect 5534 5108 5540 5160
rect 5592 5148 5598 5160
rect 5701 5151 5759 5157
rect 5701 5148 5713 5151
rect 5592 5120 5713 5148
rect 5592 5108 5598 5120
rect 5701 5117 5713 5120
rect 5747 5117 5759 5151
rect 5701 5111 5759 5117
rect 7190 5108 7196 5160
rect 7248 5108 7254 5160
rect 7285 5151 7343 5157
rect 7285 5117 7297 5151
rect 7331 5148 7343 5151
rect 7558 5148 7564 5160
rect 7331 5120 7564 5148
rect 7331 5117 7343 5120
rect 7285 5111 7343 5117
rect 7558 5108 7564 5120
rect 7616 5108 7622 5160
rect 7668 5157 7696 5256
rect 8846 5176 8852 5228
rect 8904 5216 8910 5228
rect 9493 5219 9551 5225
rect 9493 5216 9505 5219
rect 8904 5188 9505 5216
rect 8904 5176 8910 5188
rect 9493 5185 9505 5188
rect 9539 5185 9551 5219
rect 9493 5179 9551 5185
rect 12986 5176 12992 5228
rect 13044 5216 13050 5228
rect 13044 5188 13216 5216
rect 13044 5176 13050 5188
rect 7653 5151 7711 5157
rect 7653 5117 7665 5151
rect 7699 5148 7711 5151
rect 9398 5148 9404 5160
rect 7699 5120 9404 5148
rect 7699 5117 7711 5120
rect 7653 5111 7711 5117
rect 9398 5108 9404 5120
rect 9456 5108 9462 5160
rect 12066 5108 12072 5160
rect 12124 5157 12130 5160
rect 12124 5148 12136 5157
rect 12345 5151 12403 5157
rect 12124 5120 12169 5148
rect 12124 5111 12136 5120
rect 12345 5117 12357 5151
rect 12391 5117 12403 5151
rect 12345 5111 12403 5117
rect 12124 5108 12130 5111
rect 3326 5040 3332 5092
rect 3384 5040 3390 5092
rect 6454 5040 6460 5092
rect 6512 5080 6518 5092
rect 8018 5080 8024 5092
rect 6512 5052 8024 5080
rect 6512 5040 6518 5052
rect 8018 5040 8024 5052
rect 8076 5040 8082 5092
rect 8570 5040 8576 5092
rect 8628 5040 8634 5092
rect 8789 5083 8847 5089
rect 8789 5049 8801 5083
rect 8835 5080 8847 5083
rect 9033 5083 9091 5089
rect 9033 5080 9045 5083
rect 8835 5052 9045 5080
rect 8835 5049 8847 5052
rect 8789 5043 8847 5049
rect 9033 5049 9045 5052
rect 9079 5049 9091 5083
rect 9033 5043 9091 5049
rect 9217 5083 9275 5089
rect 9217 5049 9229 5083
rect 9263 5049 9275 5083
rect 9217 5043 9275 5049
rect 9760 5083 9818 5089
rect 9760 5049 9772 5083
rect 9806 5080 9818 5083
rect 10134 5080 10140 5092
rect 9806 5052 10140 5080
rect 9806 5049 9818 5052
rect 9760 5043 9818 5049
rect 2498 4972 2504 5024
rect 2556 4972 2562 5024
rect 2685 5015 2743 5021
rect 2685 4981 2697 5015
rect 2731 5012 2743 5015
rect 3234 5012 3240 5024
rect 2731 4984 3240 5012
rect 2731 4981 2743 4984
rect 2685 4975 2743 4981
rect 3234 4972 3240 4984
rect 3292 4972 3298 5024
rect 3418 4972 3424 5024
rect 3476 5012 3482 5024
rect 3529 5015 3587 5021
rect 3529 5012 3541 5015
rect 3476 4984 3541 5012
rect 3476 4972 3482 4984
rect 3529 4981 3541 4984
rect 3575 4981 3587 5015
rect 3529 4975 3587 4981
rect 3694 4972 3700 5024
rect 3752 4972 3758 5024
rect 7374 4972 7380 5024
rect 7432 4972 7438 5024
rect 8938 4972 8944 5024
rect 8996 4972 9002 5024
rect 9232 5012 9260 5043
rect 10134 5040 10140 5052
rect 10192 5040 10198 5092
rect 11422 5040 11428 5092
rect 11480 5080 11486 5092
rect 12360 5080 12388 5111
rect 12894 5108 12900 5160
rect 12952 5148 12958 5160
rect 13188 5157 13216 5188
rect 16482 5176 16488 5228
rect 16540 5176 16546 5228
rect 19168 5216 19196 5312
rect 19337 5287 19395 5293
rect 19337 5253 19349 5287
rect 19383 5284 19395 5287
rect 19794 5284 19800 5296
rect 19383 5256 19800 5284
rect 19383 5253 19395 5256
rect 19337 5247 19395 5253
rect 19794 5244 19800 5256
rect 19852 5244 19858 5296
rect 19168 5188 20576 5216
rect 13173 5151 13231 5157
rect 12952 5120 13124 5148
rect 12952 5108 12958 5120
rect 11480 5052 12388 5080
rect 11480 5040 11486 5052
rect 12526 5040 12532 5092
rect 12584 5040 12590 5092
rect 12745 5083 12803 5089
rect 12745 5049 12757 5083
rect 12791 5080 12803 5083
rect 12989 5083 13047 5089
rect 12989 5080 13001 5083
rect 12791 5052 13001 5080
rect 12791 5049 12803 5052
rect 12745 5043 12803 5049
rect 12989 5049 13001 5052
rect 13035 5049 13047 5083
rect 13096 5080 13124 5120
rect 13173 5117 13185 5151
rect 13219 5117 13231 5151
rect 13173 5111 13231 5117
rect 13354 5108 13360 5160
rect 13412 5108 13418 5160
rect 13814 5157 13820 5160
rect 13541 5151 13599 5157
rect 13541 5117 13553 5151
rect 13587 5117 13599 5151
rect 13808 5148 13820 5157
rect 13775 5120 13820 5148
rect 13541 5111 13599 5117
rect 13808 5111 13820 5120
rect 13556 5080 13584 5111
rect 13814 5108 13820 5111
rect 13872 5108 13878 5160
rect 15378 5108 15384 5160
rect 15436 5148 15442 5160
rect 16218 5151 16276 5157
rect 16218 5148 16230 5151
rect 15436 5120 16230 5148
rect 15436 5108 15442 5120
rect 16218 5117 16230 5120
rect 16264 5117 16276 5151
rect 16218 5111 16276 5117
rect 16500 5080 16528 5176
rect 20254 5108 20260 5160
rect 20312 5108 20318 5160
rect 20346 5108 20352 5160
rect 20404 5108 20410 5160
rect 20441 5151 20499 5157
rect 20441 5117 20453 5151
rect 20487 5117 20499 5151
rect 20548 5148 20576 5188
rect 20625 5151 20683 5157
rect 20625 5148 20637 5151
rect 20548 5120 20637 5148
rect 20441 5111 20499 5117
rect 20625 5117 20637 5120
rect 20671 5117 20683 5151
rect 20625 5111 20683 5117
rect 13096 5052 16528 5080
rect 18969 5083 19027 5089
rect 12989 5043 13047 5049
rect 18969 5049 18981 5083
rect 19015 5080 19027 5083
rect 20070 5080 20076 5092
rect 19015 5052 20076 5080
rect 19015 5049 19027 5052
rect 18969 5043 19027 5049
rect 20070 5040 20076 5052
rect 20128 5040 20134 5092
rect 10042 5012 10048 5024
rect 9232 4984 10048 5012
rect 10042 4972 10048 4984
rect 10100 4972 10106 5024
rect 12894 4972 12900 5024
rect 12952 4972 12958 5024
rect 14274 4972 14280 5024
rect 14332 5012 14338 5024
rect 14921 5015 14979 5021
rect 14921 5012 14933 5015
rect 14332 4984 14933 5012
rect 14332 4972 14338 4984
rect 14921 4981 14933 4984
rect 14967 4981 14979 5015
rect 14921 4975 14979 4981
rect 19978 4972 19984 5024
rect 20036 4972 20042 5024
rect 20456 5012 20484 5111
rect 20714 5108 20720 5160
rect 20772 5108 20778 5160
rect 20898 5108 20904 5160
rect 20956 5108 20962 5160
rect 21913 5151 21971 5157
rect 21913 5117 21925 5151
rect 21959 5148 21971 5151
rect 22186 5148 22192 5160
rect 21959 5120 22192 5148
rect 21959 5117 21971 5120
rect 21913 5111 21971 5117
rect 22186 5108 22192 5120
rect 22244 5108 22250 5160
rect 20809 5015 20867 5021
rect 20809 5012 20821 5015
rect 20456 4984 20821 5012
rect 20809 4981 20821 4984
rect 20855 4981 20867 5015
rect 20809 4975 20867 4981
rect 552 4922 23368 4944
rect 552 4870 4322 4922
rect 4374 4870 4386 4922
rect 4438 4870 4450 4922
rect 4502 4870 4514 4922
rect 4566 4870 4578 4922
rect 4630 4870 23368 4922
rect 552 4848 23368 4870
rect 3789 4811 3847 4817
rect 3789 4777 3801 4811
rect 3835 4808 3847 4811
rect 4062 4808 4068 4820
rect 3835 4780 4068 4808
rect 3835 4777 3847 4780
rect 3789 4771 3847 4777
rect 4062 4768 4068 4780
rect 4120 4808 4126 4820
rect 4157 4811 4215 4817
rect 4157 4808 4169 4811
rect 4120 4780 4169 4808
rect 4120 4768 4126 4780
rect 4157 4777 4169 4780
rect 4203 4777 4215 4811
rect 4157 4771 4215 4777
rect 6546 4768 6552 4820
rect 6604 4768 6610 4820
rect 8018 4768 8024 4820
rect 8076 4768 8082 4820
rect 8570 4808 8576 4820
rect 8128 4780 8576 4808
rect 2498 4700 2504 4752
rect 2556 4740 2562 4752
rect 2654 4743 2712 4749
rect 2654 4740 2666 4743
rect 2556 4712 2666 4740
rect 2556 4700 2562 4712
rect 2654 4709 2666 4712
rect 2700 4709 2712 4743
rect 2654 4703 2712 4709
rect 2866 4700 2872 4752
rect 2924 4700 2930 4752
rect 3878 4700 3884 4752
rect 3936 4700 3942 4752
rect 4706 4749 4712 4752
rect 4693 4743 4712 4749
rect 4693 4709 4705 4743
rect 4693 4703 4712 4709
rect 4706 4700 4712 4703
rect 4764 4700 4770 4752
rect 4893 4743 4951 4749
rect 4893 4709 4905 4743
rect 4939 4740 4951 4743
rect 5626 4740 5632 4752
rect 4939 4712 5632 4740
rect 4939 4709 4951 4712
rect 4893 4703 4951 4709
rect 5626 4700 5632 4712
rect 5684 4700 5690 4752
rect 5718 4700 5724 4752
rect 5776 4740 5782 4752
rect 6181 4743 6239 4749
rect 6181 4740 6193 4743
rect 5776 4712 6193 4740
rect 5776 4700 5782 4712
rect 6181 4709 6193 4712
rect 6227 4709 6239 4743
rect 6181 4703 6239 4709
rect 6717 4743 6775 4749
rect 6717 4709 6729 4743
rect 6763 4740 6775 4743
rect 6763 4709 6776 4740
rect 6717 4703 6776 4709
rect 1670 4632 1676 4684
rect 1728 4672 1734 4684
rect 2409 4675 2467 4681
rect 2409 4672 2421 4675
rect 1728 4644 2421 4672
rect 1728 4632 1734 4644
rect 2409 4641 2421 4644
rect 2455 4672 2467 4675
rect 2884 4672 2912 4700
rect 3050 4672 3056 4684
rect 2455 4644 3056 4672
rect 2455 4641 2467 4644
rect 2409 4635 2467 4641
rect 3050 4632 3056 4644
rect 3108 4632 3114 4684
rect 3142 4632 3148 4684
rect 3200 4672 3206 4684
rect 4065 4675 4123 4681
rect 4065 4672 4077 4675
rect 3200 4644 4077 4672
rect 3200 4632 3206 4644
rect 4065 4641 4077 4644
rect 4111 4641 4123 4675
rect 4065 4635 4123 4641
rect 4154 4632 4160 4684
rect 4212 4672 4218 4684
rect 4249 4675 4307 4681
rect 4249 4672 4261 4675
rect 4212 4644 4261 4672
rect 4212 4632 4218 4644
rect 4249 4641 4261 4644
rect 4295 4641 4307 4675
rect 4249 4635 4307 4641
rect 6365 4675 6423 4681
rect 6365 4641 6377 4675
rect 6411 4641 6423 4675
rect 6365 4635 6423 4641
rect 2314 4564 2320 4616
rect 2372 4564 2378 4616
rect 4264 4576 4752 4604
rect 2041 4539 2099 4545
rect 2041 4505 2053 4539
rect 2087 4505 2099 4539
rect 2041 4499 2099 4505
rect 1762 4428 1768 4480
rect 1820 4468 1826 4480
rect 1857 4471 1915 4477
rect 1857 4468 1869 4471
rect 1820 4440 1869 4468
rect 1820 4428 1826 4440
rect 1857 4437 1869 4440
rect 1903 4437 1915 4471
rect 2056 4468 2084 4499
rect 2774 4468 2780 4480
rect 2056 4440 2780 4468
rect 1857 4431 1915 4437
rect 2774 4428 2780 4440
rect 2832 4468 2838 4480
rect 4264 4468 4292 4576
rect 4430 4496 4436 4548
rect 4488 4496 4494 4548
rect 2832 4440 4292 4468
rect 2832 4428 2838 4440
rect 4338 4428 4344 4480
rect 4396 4468 4402 4480
rect 4724 4477 4752 4576
rect 6380 4536 6408 4635
rect 6748 4604 6776 4703
rect 6822 4700 6828 4752
rect 6880 4740 6886 4752
rect 8128 4749 8156 4780
rect 8570 4768 8576 4780
rect 8628 4808 8634 4820
rect 8628 4780 9076 4808
rect 8628 4768 8634 4780
rect 8938 4749 8944 4752
rect 6917 4743 6975 4749
rect 6917 4740 6929 4743
rect 6880 4712 6929 4740
rect 6880 4700 6886 4712
rect 6917 4709 6929 4712
rect 6963 4709 6975 4743
rect 6917 4703 6975 4709
rect 8113 4743 8171 4749
rect 8113 4709 8125 4743
rect 8159 4709 8171 4743
rect 8932 4740 8944 4749
rect 8899 4712 8944 4740
rect 8113 4703 8171 4709
rect 8932 4703 8944 4712
rect 8938 4700 8944 4703
rect 8996 4700 9002 4752
rect 9048 4740 9076 4780
rect 10134 4768 10140 4820
rect 10192 4768 10198 4820
rect 10321 4811 10379 4817
rect 10321 4777 10333 4811
rect 10367 4808 10379 4811
rect 11882 4808 11888 4820
rect 10367 4780 11888 4808
rect 10367 4777 10379 4780
rect 10321 4771 10379 4777
rect 10336 4740 10364 4771
rect 11882 4768 11888 4780
rect 11940 4768 11946 4820
rect 13722 4768 13728 4820
rect 13780 4808 13786 4820
rect 14185 4811 14243 4817
rect 14185 4808 14197 4811
rect 13780 4780 14197 4808
rect 13780 4768 13786 4780
rect 14185 4777 14197 4780
rect 14231 4777 14243 4811
rect 14185 4771 14243 4777
rect 20254 4768 20260 4820
rect 20312 4808 20318 4820
rect 20898 4808 20904 4820
rect 20312 4780 20904 4808
rect 20312 4768 20318 4780
rect 20898 4768 20904 4780
rect 20956 4808 20962 4820
rect 21085 4811 21143 4817
rect 21085 4808 21097 4811
rect 20956 4780 21097 4808
rect 20956 4768 20962 4780
rect 21085 4777 21097 4780
rect 21131 4777 21143 4811
rect 21085 4771 21143 4777
rect 9048 4712 10364 4740
rect 12894 4700 12900 4752
rect 12952 4740 12958 4752
rect 19978 4749 19984 4752
rect 13050 4743 13108 4749
rect 13050 4740 13062 4743
rect 12952 4712 13062 4740
rect 12952 4700 12958 4712
rect 13050 4709 13062 4712
rect 13096 4709 13108 4743
rect 19972 4740 19984 4749
rect 19939 4712 19984 4740
rect 13050 4703 13108 4709
rect 19972 4703 19984 4712
rect 19978 4700 19984 4703
rect 20036 4700 20042 4752
rect 8754 4672 8760 4684
rect 8680 4644 8760 4672
rect 7374 4604 7380 4616
rect 6748 4576 7380 4604
rect 7374 4564 7380 4576
rect 7432 4564 7438 4616
rect 8680 4613 8708 4644
rect 8754 4632 8760 4644
rect 8812 4632 8818 4684
rect 11422 4632 11428 4684
rect 11480 4672 11486 4684
rect 11517 4675 11575 4681
rect 11517 4672 11529 4675
rect 11480 4644 11529 4672
rect 11480 4632 11486 4644
rect 11517 4641 11529 4644
rect 11563 4641 11575 4675
rect 11517 4635 11575 4641
rect 11793 4675 11851 4681
rect 11793 4641 11805 4675
rect 11839 4672 11851 4675
rect 11839 4644 22094 4672
rect 11839 4641 11851 4644
rect 11793 4635 11851 4641
rect 8665 4607 8723 4613
rect 8665 4573 8677 4607
rect 8711 4573 8723 4607
rect 8665 4567 8723 4573
rect 8680 4536 8708 4567
rect 12802 4564 12808 4616
rect 12860 4564 12866 4616
rect 19702 4564 19708 4616
rect 19760 4564 19766 4616
rect 6380 4508 8708 4536
rect 10226 4496 10232 4548
rect 10284 4536 10290 4548
rect 10689 4539 10747 4545
rect 10689 4536 10701 4539
rect 10284 4508 10701 4536
rect 10284 4496 10290 4508
rect 10689 4505 10701 4508
rect 10735 4505 10747 4539
rect 10689 4499 10747 4505
rect 4525 4471 4583 4477
rect 4525 4468 4537 4471
rect 4396 4440 4537 4468
rect 4396 4428 4402 4440
rect 4525 4437 4537 4440
rect 4571 4437 4583 4471
rect 4525 4431 4583 4437
rect 4709 4471 4767 4477
rect 4709 4437 4721 4471
rect 4755 4437 4767 4471
rect 4709 4431 4767 4437
rect 6733 4471 6791 4477
rect 6733 4437 6745 4471
rect 6779 4468 6791 4471
rect 7190 4468 7196 4480
rect 6779 4440 7196 4468
rect 6779 4437 6791 4440
rect 6733 4431 6791 4437
rect 7190 4428 7196 4440
rect 7248 4428 7254 4480
rect 10042 4428 10048 4480
rect 10100 4428 10106 4480
rect 10318 4428 10324 4480
rect 10376 4428 10382 4480
rect 22066 4468 22094 4644
rect 22462 4468 22468 4480
rect 22066 4440 22468 4468
rect 22462 4428 22468 4440
rect 22520 4468 22526 4480
rect 22830 4468 22836 4480
rect 22520 4440 22836 4468
rect 22520 4428 22526 4440
rect 22830 4428 22836 4440
rect 22888 4428 22894 4480
rect 552 4378 23368 4400
rect 552 4326 3662 4378
rect 3714 4326 3726 4378
rect 3778 4326 3790 4378
rect 3842 4326 3854 4378
rect 3906 4326 3918 4378
rect 3970 4326 23368 4378
rect 552 4304 23368 4326
rect 2314 4224 2320 4276
rect 2372 4264 2378 4276
rect 2866 4264 2872 4276
rect 2372 4236 2872 4264
rect 2372 4224 2378 4236
rect 2866 4224 2872 4236
rect 2924 4264 2930 4276
rect 3053 4267 3111 4273
rect 3053 4264 3065 4267
rect 2924 4236 3065 4264
rect 2924 4224 2930 4236
rect 3053 4233 3065 4236
rect 3099 4233 3111 4267
rect 4430 4264 4436 4276
rect 3053 4227 3111 4233
rect 3620 4236 4436 4264
rect 3068 4196 3096 4227
rect 3620 4196 3648 4236
rect 4430 4224 4436 4236
rect 4488 4264 4494 4276
rect 4798 4264 4804 4276
rect 4488 4236 4804 4264
rect 4488 4224 4494 4236
rect 4798 4224 4804 4236
rect 4856 4224 4862 4276
rect 10226 4224 10232 4276
rect 10284 4224 10290 4276
rect 10413 4267 10471 4273
rect 10413 4233 10425 4267
rect 10459 4264 10471 4267
rect 10686 4264 10692 4276
rect 10459 4236 10692 4264
rect 10459 4233 10471 4236
rect 10413 4227 10471 4233
rect 10686 4224 10692 4236
rect 10744 4224 10750 4276
rect 22830 4224 22836 4276
rect 22888 4224 22894 4276
rect 3068 4168 3648 4196
rect 1670 4088 1676 4140
rect 1728 4088 1734 4140
rect 3234 4088 3240 4140
rect 3292 4088 3298 4140
rect 3620 4137 3648 4168
rect 4062 4156 4068 4208
rect 4120 4156 4126 4208
rect 3605 4131 3663 4137
rect 3605 4097 3617 4131
rect 3651 4097 3663 4131
rect 3605 4091 3663 4097
rect 3697 4131 3755 4137
rect 3697 4097 3709 4131
rect 3743 4128 3755 4131
rect 4080 4128 4108 4156
rect 3743 4100 4108 4128
rect 3743 4097 3755 4100
rect 3697 4091 3755 4097
rect 5626 4088 5632 4140
rect 5684 4088 5690 4140
rect 11333 4131 11391 4137
rect 11333 4097 11345 4131
rect 11379 4128 11391 4131
rect 11974 4128 11980 4140
rect 11379 4100 11980 4128
rect 11379 4097 11391 4100
rect 11333 4091 11391 4097
rect 11974 4088 11980 4100
rect 12032 4088 12038 4140
rect 1762 4020 1768 4072
rect 1820 4060 1826 4072
rect 1929 4063 1987 4069
rect 1929 4060 1941 4063
rect 1820 4032 1941 4060
rect 1820 4020 1826 4032
rect 1929 4029 1941 4032
rect 1975 4029 1987 4063
rect 1929 4023 1987 4029
rect 3142 4020 3148 4072
rect 3200 4060 3206 4072
rect 3421 4063 3479 4069
rect 3421 4060 3433 4063
rect 3200 4032 3433 4060
rect 3200 4020 3206 4032
rect 3421 4029 3433 4032
rect 3467 4029 3479 4063
rect 3421 4023 3479 4029
rect 3513 4063 3571 4069
rect 3513 4029 3525 4063
rect 3559 4029 3571 4063
rect 3513 4023 3571 4029
rect 2958 3952 2964 4004
rect 3016 3992 3022 4004
rect 3528 3992 3556 4023
rect 4062 4020 4068 4072
rect 4120 4020 4126 4072
rect 4338 4069 4344 4072
rect 4332 4060 4344 4069
rect 4299 4032 4344 4060
rect 4332 4023 4344 4032
rect 4338 4020 4344 4023
rect 4396 4020 4402 4072
rect 4798 4020 4804 4072
rect 4856 4060 4862 4072
rect 5537 4063 5595 4069
rect 5537 4060 5549 4063
rect 4856 4032 5549 4060
rect 4856 4020 4862 4032
rect 5537 4029 5549 4032
rect 5583 4029 5595 4063
rect 5537 4023 5595 4029
rect 5721 4063 5779 4069
rect 5721 4029 5733 4063
rect 5767 4029 5779 4063
rect 5721 4023 5779 4029
rect 4154 3992 4160 4004
rect 3016 3964 4160 3992
rect 3016 3952 3022 3964
rect 4154 3952 4160 3964
rect 4212 3952 4218 4004
rect 5736 3992 5764 4023
rect 10226 4020 10232 4072
rect 10284 4060 10290 4072
rect 10965 4063 11023 4069
rect 10965 4060 10977 4063
rect 10284 4032 10977 4060
rect 10284 4020 10290 4032
rect 10965 4029 10977 4032
rect 11011 4029 11023 4063
rect 10965 4023 11023 4029
rect 11146 4020 11152 4072
rect 11204 4020 11210 4072
rect 23014 4020 23020 4072
rect 23072 4020 23078 4072
rect 5460 3964 5764 3992
rect 5460 3936 5488 3964
rect 10042 3952 10048 4004
rect 10100 3992 10106 4004
rect 10597 3995 10655 4001
rect 10597 3992 10609 3995
rect 10100 3964 10609 3992
rect 10100 3952 10106 3964
rect 10597 3961 10609 3964
rect 10643 3961 10655 3995
rect 10597 3955 10655 3961
rect 5442 3884 5448 3936
rect 5500 3884 5506 3936
rect 9398 3884 9404 3936
rect 9456 3924 9462 3936
rect 10387 3927 10445 3933
rect 10387 3924 10399 3927
rect 9456 3896 10399 3924
rect 9456 3884 9462 3896
rect 10387 3893 10399 3896
rect 10433 3893 10445 3927
rect 10387 3887 10445 3893
rect 552 3834 23368 3856
rect 552 3782 4322 3834
rect 4374 3782 4386 3834
rect 4438 3782 4450 3834
rect 4502 3782 4514 3834
rect 4566 3782 4578 3834
rect 4630 3782 23368 3834
rect 552 3760 23368 3782
rect 3053 3723 3111 3729
rect 3053 3689 3065 3723
rect 3099 3720 3111 3723
rect 3326 3720 3332 3732
rect 3099 3692 3332 3720
rect 3099 3689 3111 3692
rect 3053 3683 3111 3689
rect 3326 3680 3332 3692
rect 3384 3680 3390 3732
rect 4617 3723 4675 3729
rect 4617 3720 4629 3723
rect 3420 3692 4629 3720
rect 2958 3612 2964 3664
rect 3016 3612 3022 3664
rect 3142 3612 3148 3664
rect 3200 3652 3206 3664
rect 3420 3652 3448 3692
rect 4617 3689 4629 3692
rect 4663 3689 4675 3723
rect 4617 3683 4675 3689
rect 4706 3680 4712 3732
rect 4764 3680 4770 3732
rect 3510 3661 3516 3664
rect 3200 3624 3448 3652
rect 3200 3612 3206 3624
rect 3504 3615 3516 3661
rect 3568 3652 3574 3664
rect 3568 3624 3604 3652
rect 3510 3612 3516 3615
rect 3568 3612 3574 3624
rect 4154 3612 4160 3664
rect 4212 3652 4218 3664
rect 5077 3655 5135 3661
rect 5077 3652 5089 3655
rect 4212 3624 5089 3652
rect 4212 3612 4218 3624
rect 5077 3621 5089 3624
rect 5123 3652 5135 3655
rect 5442 3652 5448 3664
rect 5123 3624 5448 3652
rect 5123 3621 5135 3624
rect 5077 3615 5135 3621
rect 5442 3612 5448 3624
rect 5500 3612 5506 3664
rect 2866 3544 2872 3596
rect 2924 3544 2930 3596
rect 3050 3544 3056 3596
rect 3108 3584 3114 3596
rect 3237 3587 3295 3593
rect 3237 3584 3249 3587
rect 3108 3556 3249 3584
rect 3108 3544 3114 3556
rect 3237 3553 3249 3556
rect 3283 3584 3295 3587
rect 4062 3584 4068 3596
rect 3283 3556 4068 3584
rect 3283 3553 3295 3556
rect 3237 3547 3295 3553
rect 4062 3544 4068 3556
rect 4120 3544 4126 3596
rect 4798 3544 4804 3596
rect 4856 3584 4862 3596
rect 4893 3587 4951 3593
rect 4893 3584 4905 3587
rect 4856 3556 4905 3584
rect 4856 3544 4862 3556
rect 4893 3553 4905 3556
rect 4939 3553 4951 3587
rect 4893 3547 4951 3553
rect 552 3290 23368 3312
rect 552 3238 3662 3290
rect 3714 3238 3726 3290
rect 3778 3238 3790 3290
rect 3842 3238 3854 3290
rect 3906 3238 3918 3290
rect 3970 3238 23368 3290
rect 552 3216 23368 3238
rect 3418 3136 3424 3188
rect 3476 3136 3482 3188
rect 2866 3000 2872 3052
rect 2924 3040 2930 3052
rect 2924 3012 3832 3040
rect 2924 3000 2930 3012
rect 3142 2932 3148 2984
rect 3200 2972 3206 2984
rect 3804 2981 3832 3012
rect 3605 2975 3663 2981
rect 3605 2972 3617 2975
rect 3200 2944 3617 2972
rect 3200 2932 3206 2944
rect 3605 2941 3617 2944
rect 3651 2941 3663 2975
rect 3605 2935 3663 2941
rect 3789 2975 3847 2981
rect 3789 2941 3801 2975
rect 3835 2941 3847 2975
rect 3789 2935 3847 2941
rect 3881 2975 3939 2981
rect 3881 2941 3893 2975
rect 3927 2972 3939 2975
rect 4154 2972 4160 2984
rect 3927 2944 4160 2972
rect 3927 2941 3939 2944
rect 3881 2935 3939 2941
rect 4154 2932 4160 2944
rect 4212 2932 4218 2984
rect 552 2746 23368 2768
rect 552 2694 4322 2746
rect 4374 2694 4386 2746
rect 4438 2694 4450 2746
rect 4502 2694 4514 2746
rect 4566 2694 4578 2746
rect 4630 2694 23368 2746
rect 552 2672 23368 2694
rect 552 2202 23368 2224
rect 552 2150 3662 2202
rect 3714 2150 3726 2202
rect 3778 2150 3790 2202
rect 3842 2150 3854 2202
rect 3906 2150 3918 2202
rect 3970 2150 23368 2202
rect 552 2128 23368 2150
rect 552 1658 23368 1680
rect 552 1606 4322 1658
rect 4374 1606 4386 1658
rect 4438 1606 4450 1658
rect 4502 1606 4514 1658
rect 4566 1606 4578 1658
rect 4630 1606 23368 1658
rect 552 1584 23368 1606
rect 552 1114 23368 1136
rect 552 1062 3662 1114
rect 3714 1062 3726 1114
rect 3778 1062 3790 1114
rect 3842 1062 3854 1114
rect 3906 1062 3918 1114
rect 3970 1062 23368 1114
rect 552 1040 23368 1062
rect 552 570 23368 592
rect 552 518 4322 570
rect 4374 518 4386 570
rect 4438 518 4450 570
rect 4502 518 4514 570
rect 4566 518 4578 570
rect 4630 518 23368 570
rect 552 496 23368 518
<< via1 >>
rect 4322 23366 4374 23418
rect 4386 23366 4438 23418
rect 4450 23366 4502 23418
rect 4514 23366 4566 23418
rect 4578 23366 4630 23418
rect 5264 23264 5316 23316
rect 3424 23196 3476 23248
rect 1768 23171 1820 23180
rect 1768 23137 1777 23171
rect 1777 23137 1811 23171
rect 1811 23137 1820 23171
rect 1768 23128 1820 23137
rect 2780 23128 2832 23180
rect 4896 23196 4948 23248
rect 3424 23060 3476 23112
rect 4344 23128 4396 23180
rect 4988 23171 5040 23180
rect 4988 23137 4997 23171
rect 4997 23137 5031 23171
rect 5031 23137 5040 23171
rect 4988 23128 5040 23137
rect 5264 23128 5316 23180
rect 10508 23196 10560 23248
rect 7564 23128 7616 23180
rect 13544 23171 13596 23180
rect 13544 23137 13553 23171
rect 13553 23137 13587 23171
rect 13587 23137 13596 23171
rect 13544 23128 13596 23137
rect 16488 23171 16540 23180
rect 16488 23137 16497 23171
rect 16497 23137 16531 23171
rect 16531 23137 16540 23171
rect 16488 23128 16540 23137
rect 17960 23128 18012 23180
rect 18788 23128 18840 23180
rect 19432 23171 19484 23180
rect 19432 23137 19441 23171
rect 19441 23137 19475 23171
rect 19475 23137 19484 23171
rect 19432 23128 19484 23137
rect 22284 23128 22336 23180
rect 5816 23060 5868 23112
rect 13912 23060 13964 23112
rect 15200 23060 15252 23112
rect 15476 23060 15528 23112
rect 18420 23060 18472 23112
rect 21916 23060 21968 23112
rect 22008 23060 22060 23112
rect 2872 22992 2924 23044
rect 3056 22924 3108 22976
rect 7288 22992 7340 23044
rect 21456 22992 21508 23044
rect 7196 22924 7248 22976
rect 9588 22924 9640 22976
rect 14096 22924 14148 22976
rect 16672 22967 16724 22976
rect 16672 22933 16681 22967
rect 16681 22933 16715 22967
rect 16715 22933 16724 22967
rect 16672 22924 16724 22933
rect 18328 22967 18380 22976
rect 18328 22933 18337 22967
rect 18337 22933 18371 22967
rect 18371 22933 18380 22967
rect 18328 22924 18380 22933
rect 3662 22822 3714 22874
rect 3726 22822 3778 22874
rect 3790 22822 3842 22874
rect 3854 22822 3906 22874
rect 3918 22822 3970 22874
rect 4712 22720 4764 22772
rect 7196 22720 7248 22772
rect 7288 22720 7340 22772
rect 8208 22720 8260 22772
rect 6000 22652 6052 22704
rect 3056 22559 3108 22568
rect 3056 22525 3065 22559
rect 3065 22525 3099 22559
rect 3099 22525 3108 22559
rect 3056 22516 3108 22525
rect 3424 22559 3476 22568
rect 3424 22525 3433 22559
rect 3433 22525 3467 22559
rect 3467 22525 3476 22559
rect 3424 22516 3476 22525
rect 14004 22720 14056 22772
rect 15292 22720 15344 22772
rect 4344 22516 4396 22568
rect 4712 22559 4764 22568
rect 4712 22525 4721 22559
rect 4721 22525 4755 22559
rect 4755 22525 4764 22559
rect 4712 22516 4764 22525
rect 4804 22516 4856 22568
rect 6276 22516 6328 22568
rect 7472 22516 7524 22568
rect 7840 22516 7892 22568
rect 8484 22516 8536 22568
rect 10600 22516 10652 22568
rect 11796 22559 11848 22568
rect 11796 22525 11805 22559
rect 11805 22525 11839 22559
rect 11839 22525 11848 22559
rect 11796 22516 11848 22525
rect 12532 22559 12584 22568
rect 12532 22525 12541 22559
rect 12541 22525 12575 22559
rect 12575 22525 12584 22559
rect 12532 22516 12584 22525
rect 13820 22584 13872 22636
rect 5080 22448 5132 22500
rect 7748 22448 7800 22500
rect 2872 22423 2924 22432
rect 2872 22389 2881 22423
rect 2881 22389 2915 22423
rect 2915 22389 2924 22423
rect 2872 22380 2924 22389
rect 7104 22380 7156 22432
rect 7932 22380 7984 22432
rect 8208 22380 8260 22432
rect 10416 22448 10468 22500
rect 12072 22491 12124 22500
rect 12072 22457 12081 22491
rect 12081 22457 12115 22491
rect 12115 22457 12124 22491
rect 12072 22448 12124 22457
rect 12440 22448 12492 22500
rect 12808 22559 12860 22568
rect 12808 22525 12818 22559
rect 12818 22525 12852 22559
rect 12852 22525 12860 22559
rect 12808 22516 12860 22525
rect 12900 22448 12952 22500
rect 8668 22380 8720 22432
rect 10324 22423 10376 22432
rect 10324 22389 10333 22423
rect 10333 22389 10367 22423
rect 10367 22389 10376 22423
rect 10324 22380 10376 22389
rect 11704 22380 11756 22432
rect 12256 22423 12308 22432
rect 12256 22389 12265 22423
rect 12265 22389 12299 22423
rect 12299 22389 12308 22423
rect 12256 22380 12308 22389
rect 12716 22380 12768 22432
rect 17960 22720 18012 22772
rect 14096 22559 14148 22568
rect 14096 22525 14105 22559
rect 14105 22525 14139 22559
rect 14139 22525 14148 22559
rect 14096 22516 14148 22525
rect 14188 22448 14240 22500
rect 15292 22516 15344 22568
rect 15200 22491 15252 22500
rect 15200 22457 15209 22491
rect 15209 22457 15243 22491
rect 15243 22457 15252 22491
rect 15200 22448 15252 22457
rect 14832 22380 14884 22432
rect 15016 22423 15068 22432
rect 15016 22389 15025 22423
rect 15025 22389 15059 22423
rect 15059 22389 15068 22423
rect 15016 22380 15068 22389
rect 15292 22423 15344 22432
rect 15292 22389 15301 22423
rect 15301 22389 15335 22423
rect 15335 22389 15344 22423
rect 15292 22380 15344 22389
rect 16856 22516 16908 22568
rect 18328 22584 18380 22636
rect 18420 22559 18472 22568
rect 15660 22491 15712 22500
rect 15660 22457 15669 22491
rect 15669 22457 15703 22491
rect 15703 22457 15712 22491
rect 15660 22448 15712 22457
rect 16672 22491 16724 22500
rect 16672 22457 16681 22491
rect 16681 22457 16715 22491
rect 16715 22457 16724 22491
rect 16672 22448 16724 22457
rect 18420 22525 18429 22559
rect 18429 22525 18463 22559
rect 18463 22525 18472 22559
rect 18420 22516 18472 22525
rect 19248 22516 19300 22568
rect 20076 22516 20128 22568
rect 20720 22584 20772 22636
rect 21364 22627 21416 22636
rect 21364 22593 21373 22627
rect 21373 22593 21407 22627
rect 21407 22593 21416 22627
rect 21364 22584 21416 22593
rect 20628 22491 20680 22500
rect 20628 22457 20637 22491
rect 20637 22457 20671 22491
rect 20671 22457 20680 22491
rect 20628 22448 20680 22457
rect 20812 22448 20864 22500
rect 21824 22448 21876 22500
rect 18788 22380 18840 22432
rect 19892 22380 19944 22432
rect 21548 22423 21600 22432
rect 21548 22389 21557 22423
rect 21557 22389 21591 22423
rect 21591 22389 21600 22423
rect 21548 22380 21600 22389
rect 4322 22278 4374 22330
rect 4386 22278 4438 22330
rect 4450 22278 4502 22330
rect 4514 22278 4566 22330
rect 4578 22278 4630 22330
rect 6276 22151 6328 22160
rect 6276 22117 6285 22151
rect 6285 22117 6319 22151
rect 6319 22117 6328 22151
rect 6276 22108 6328 22117
rect 4252 22083 4304 22092
rect 4252 22049 4261 22083
rect 4261 22049 4295 22083
rect 4295 22049 4304 22083
rect 4252 22040 4304 22049
rect 5080 22083 5132 22092
rect 5080 22049 5089 22083
rect 5089 22049 5123 22083
rect 5123 22049 5132 22083
rect 5080 22040 5132 22049
rect 5816 22083 5868 22092
rect 5816 22049 5825 22083
rect 5825 22049 5859 22083
rect 5859 22049 5868 22083
rect 5816 22040 5868 22049
rect 6000 22083 6052 22092
rect 6000 22049 6009 22083
rect 6009 22049 6043 22083
rect 6043 22049 6052 22083
rect 6828 22176 6880 22228
rect 8484 22176 8536 22228
rect 12532 22176 12584 22228
rect 13360 22219 13412 22228
rect 13360 22185 13369 22219
rect 13369 22185 13403 22219
rect 13403 22185 13412 22219
rect 13360 22176 13412 22185
rect 13912 22176 13964 22228
rect 14096 22176 14148 22228
rect 15016 22176 15068 22228
rect 8116 22108 8168 22160
rect 6000 22040 6052 22049
rect 7012 22083 7064 22092
rect 7012 22049 7021 22083
rect 7021 22049 7055 22083
rect 7055 22049 7064 22083
rect 7012 22040 7064 22049
rect 7104 22083 7156 22092
rect 7104 22049 7113 22083
rect 7113 22049 7147 22083
rect 7147 22049 7156 22083
rect 7104 22040 7156 22049
rect 7748 22083 7800 22092
rect 7748 22049 7757 22083
rect 7757 22049 7791 22083
rect 7791 22049 7800 22083
rect 7748 22040 7800 22049
rect 7932 22040 7984 22092
rect 8300 22083 8352 22092
rect 8300 22049 8309 22083
rect 8309 22049 8343 22083
rect 8343 22049 8352 22083
rect 8300 22040 8352 22049
rect 8576 22083 8628 22092
rect 8576 22049 8585 22083
rect 8585 22049 8619 22083
rect 8619 22049 8628 22083
rect 8576 22040 8628 22049
rect 8668 22083 8720 22092
rect 8668 22049 8677 22083
rect 8677 22049 8711 22083
rect 8711 22049 8720 22083
rect 8668 22040 8720 22049
rect 9312 22083 9364 22092
rect 9312 22049 9321 22083
rect 9321 22049 9355 22083
rect 9355 22049 9364 22083
rect 9312 22040 9364 22049
rect 9496 22083 9548 22092
rect 9496 22049 9505 22083
rect 9505 22049 9539 22083
rect 9539 22049 9548 22083
rect 9496 22040 9548 22049
rect 5172 21947 5224 21956
rect 5172 21913 5181 21947
rect 5181 21913 5215 21947
rect 5215 21913 5224 21947
rect 5172 21904 5224 21913
rect 6920 21972 6972 22024
rect 11796 22108 11848 22160
rect 13728 22151 13780 22160
rect 13728 22117 13737 22151
rect 13737 22117 13771 22151
rect 13771 22117 13780 22151
rect 13728 22108 13780 22117
rect 14740 22108 14792 22160
rect 15476 22151 15528 22160
rect 15476 22117 15501 22151
rect 15501 22117 15528 22151
rect 15660 22219 15712 22228
rect 15660 22185 15669 22219
rect 15669 22185 15703 22219
rect 15703 22185 15712 22219
rect 15660 22176 15712 22185
rect 16948 22176 17000 22228
rect 20628 22176 20680 22228
rect 21364 22176 21416 22228
rect 22008 22176 22060 22228
rect 15476 22108 15528 22117
rect 10416 22083 10468 22092
rect 10416 22049 10425 22083
rect 10425 22049 10459 22083
rect 10459 22049 10468 22083
rect 10416 22040 10468 22049
rect 10508 22083 10560 22092
rect 10508 22049 10518 22083
rect 10518 22049 10552 22083
rect 10552 22049 10560 22083
rect 10508 22040 10560 22049
rect 10784 22040 10836 22092
rect 10692 21972 10744 22024
rect 12808 22040 12860 22092
rect 12900 22083 12952 22092
rect 12900 22049 12909 22083
rect 12909 22049 12943 22083
rect 12943 22049 12952 22083
rect 12900 22040 12952 22049
rect 13360 22040 13412 22092
rect 13268 22015 13320 22024
rect 13268 21981 13277 22015
rect 13277 21981 13311 22015
rect 13311 21981 13320 22015
rect 13268 21972 13320 21981
rect 13820 22015 13872 22024
rect 13820 21981 13829 22015
rect 13829 21981 13863 22015
rect 13863 21981 13872 22015
rect 13820 21972 13872 21981
rect 14004 22083 14056 22092
rect 14004 22049 14013 22083
rect 14013 22049 14047 22083
rect 14047 22049 14056 22083
rect 14004 22040 14056 22049
rect 15660 22040 15712 22092
rect 16856 22083 16908 22092
rect 16856 22049 16865 22083
rect 16865 22049 16899 22083
rect 16899 22049 16908 22083
rect 16856 22040 16908 22049
rect 19248 22108 19300 22160
rect 19892 22151 19944 22160
rect 19892 22117 19901 22151
rect 19901 22117 19935 22151
rect 19935 22117 19944 22151
rect 19892 22108 19944 22117
rect 15292 21972 15344 22024
rect 16672 21972 16724 22024
rect 17960 22040 18012 22092
rect 18788 22083 18840 22092
rect 18788 22049 18797 22083
rect 18797 22049 18831 22083
rect 18831 22049 18840 22083
rect 18788 22040 18840 22049
rect 18052 21972 18104 22024
rect 18328 21972 18380 22024
rect 20352 22015 20404 22024
rect 20352 21981 20361 22015
rect 20361 21981 20395 22015
rect 20395 21981 20404 22015
rect 20352 21972 20404 21981
rect 10416 21904 10468 21956
rect 11704 21904 11756 21956
rect 5908 21879 5960 21888
rect 5908 21845 5917 21879
rect 5917 21845 5951 21879
rect 5951 21845 5960 21879
rect 5908 21836 5960 21845
rect 6368 21836 6420 21888
rect 7288 21879 7340 21888
rect 7288 21845 7297 21879
rect 7297 21845 7331 21879
rect 7331 21845 7340 21879
rect 7288 21836 7340 21845
rect 10232 21836 10284 21888
rect 14648 21947 14700 21956
rect 14648 21913 14657 21947
rect 14657 21913 14691 21947
rect 14691 21913 14700 21947
rect 14648 21904 14700 21913
rect 15016 21904 15068 21956
rect 21640 22083 21692 22092
rect 21640 22049 21649 22083
rect 21649 22049 21683 22083
rect 21683 22049 21692 22083
rect 21640 22040 21692 22049
rect 21824 22040 21876 22092
rect 22008 22074 22060 22126
rect 22100 22040 22152 22092
rect 21456 21972 21508 22024
rect 22008 21972 22060 22024
rect 20720 21904 20772 21956
rect 20996 21904 21048 21956
rect 21088 21904 21140 21956
rect 13728 21836 13780 21888
rect 14188 21836 14240 21888
rect 16304 21879 16356 21888
rect 16304 21845 16313 21879
rect 16313 21845 16347 21879
rect 16347 21845 16356 21879
rect 16304 21836 16356 21845
rect 18144 21836 18196 21888
rect 18328 21879 18380 21888
rect 18328 21845 18337 21879
rect 18337 21845 18371 21879
rect 18371 21845 18380 21879
rect 18328 21836 18380 21845
rect 19248 21836 19300 21888
rect 19524 21836 19576 21888
rect 20076 21879 20128 21888
rect 20076 21845 20085 21879
rect 20085 21845 20119 21879
rect 20119 21845 20128 21879
rect 20076 21836 20128 21845
rect 20812 21836 20864 21888
rect 20904 21879 20956 21888
rect 20904 21845 20913 21879
rect 20913 21845 20947 21879
rect 20947 21845 20956 21879
rect 20904 21836 20956 21845
rect 21180 21836 21232 21888
rect 21732 21904 21784 21956
rect 22284 22015 22336 22024
rect 22284 21981 22293 22015
rect 22293 21981 22327 22015
rect 22327 21981 22336 22015
rect 22284 21972 22336 21981
rect 22100 21879 22152 21888
rect 22100 21845 22109 21879
rect 22109 21845 22143 21879
rect 22143 21845 22152 21879
rect 22100 21836 22152 21845
rect 3662 21734 3714 21786
rect 3726 21734 3778 21786
rect 3790 21734 3842 21786
rect 3854 21734 3906 21786
rect 3918 21734 3970 21786
rect 6920 21632 6972 21684
rect 7748 21632 7800 21684
rect 8116 21632 8168 21684
rect 8576 21632 8628 21684
rect 9772 21632 9824 21684
rect 10508 21632 10560 21684
rect 12440 21632 12492 21684
rect 12900 21632 12952 21684
rect 13636 21632 13688 21684
rect 14740 21632 14792 21684
rect 15568 21632 15620 21684
rect 16764 21632 16816 21684
rect 20812 21632 20864 21684
rect 21364 21632 21416 21684
rect 21732 21632 21784 21684
rect 7564 21564 7616 21616
rect 8300 21564 8352 21616
rect 5172 21539 5224 21548
rect 5172 21505 5181 21539
rect 5181 21505 5215 21539
rect 5215 21505 5224 21539
rect 5172 21496 5224 21505
rect 6276 21496 6328 21548
rect 6828 21496 6880 21548
rect 4252 21428 4304 21480
rect 4804 21428 4856 21480
rect 5908 21428 5960 21480
rect 7472 21471 7524 21480
rect 7472 21437 7481 21471
rect 7481 21437 7515 21471
rect 7515 21437 7524 21471
rect 7472 21428 7524 21437
rect 7656 21428 7708 21480
rect 7840 21539 7892 21548
rect 7840 21505 7849 21539
rect 7849 21505 7883 21539
rect 7883 21505 7892 21539
rect 7840 21496 7892 21505
rect 8852 21564 8904 21616
rect 9496 21564 9548 21616
rect 8208 21403 8260 21412
rect 8208 21369 8220 21403
rect 8220 21369 8254 21403
rect 8254 21369 8260 21403
rect 8576 21471 8628 21480
rect 8576 21437 8585 21471
rect 8585 21437 8619 21471
rect 8619 21437 8628 21471
rect 8576 21428 8628 21437
rect 8852 21471 8904 21480
rect 8852 21437 8861 21471
rect 8861 21437 8895 21471
rect 8895 21437 8904 21471
rect 8852 21428 8904 21437
rect 8944 21471 8996 21480
rect 8944 21437 8953 21471
rect 8953 21437 8987 21471
rect 8987 21437 8996 21471
rect 8944 21428 8996 21437
rect 9220 21496 9272 21548
rect 9588 21496 9640 21548
rect 10232 21539 10284 21548
rect 10232 21505 10241 21539
rect 10241 21505 10275 21539
rect 10275 21505 10284 21539
rect 10232 21496 10284 21505
rect 8208 21360 8260 21369
rect 9036 21360 9088 21412
rect 10324 21428 10376 21480
rect 10692 21428 10744 21480
rect 12532 21564 12584 21616
rect 14096 21564 14148 21616
rect 11704 21539 11756 21548
rect 11704 21505 11713 21539
rect 11713 21505 11747 21539
rect 11747 21505 11756 21539
rect 11704 21496 11756 21505
rect 12256 21539 12308 21548
rect 12256 21505 12265 21539
rect 12265 21505 12299 21539
rect 12299 21505 12308 21539
rect 12256 21496 12308 21505
rect 12716 21539 12768 21548
rect 12716 21505 12725 21539
rect 12725 21505 12759 21539
rect 12759 21505 12768 21539
rect 12716 21496 12768 21505
rect 11796 21428 11848 21480
rect 12808 21428 12860 21480
rect 13728 21496 13780 21548
rect 9312 21360 9364 21412
rect 9404 21403 9456 21412
rect 9404 21369 9413 21403
rect 9413 21369 9447 21403
rect 9447 21369 9456 21403
rect 9404 21360 9456 21369
rect 3976 21292 4028 21344
rect 5908 21335 5960 21344
rect 5908 21301 5917 21335
rect 5917 21301 5951 21335
rect 5951 21301 5960 21335
rect 5908 21292 5960 21301
rect 6184 21292 6236 21344
rect 6368 21335 6420 21344
rect 6368 21301 6377 21335
rect 6377 21301 6411 21335
rect 6411 21301 6420 21335
rect 6368 21292 6420 21301
rect 7748 21292 7800 21344
rect 8576 21292 8628 21344
rect 8668 21292 8720 21344
rect 10140 21292 10192 21344
rect 11336 21360 11388 21412
rect 12072 21403 12124 21412
rect 12072 21369 12081 21403
rect 12081 21369 12115 21403
rect 12115 21369 12124 21403
rect 12072 21360 12124 21369
rect 12900 21360 12952 21412
rect 13268 21428 13320 21480
rect 18328 21564 18380 21616
rect 10692 21335 10744 21344
rect 10692 21301 10701 21335
rect 10701 21301 10735 21335
rect 10735 21301 10744 21335
rect 10692 21292 10744 21301
rect 11060 21335 11112 21344
rect 11060 21301 11069 21335
rect 11069 21301 11103 21335
rect 11103 21301 11112 21335
rect 11060 21292 11112 21301
rect 11152 21292 11204 21344
rect 12532 21292 12584 21344
rect 13084 21292 13136 21344
rect 13360 21335 13412 21344
rect 13360 21301 13369 21335
rect 13369 21301 13403 21335
rect 13403 21301 13412 21335
rect 13360 21292 13412 21301
rect 13544 21403 13596 21412
rect 13544 21369 13553 21403
rect 13553 21369 13587 21403
rect 13587 21369 13596 21403
rect 13544 21360 13596 21369
rect 14832 21428 14884 21480
rect 14740 21403 14792 21412
rect 14740 21369 14749 21403
rect 14749 21369 14783 21403
rect 14783 21369 14792 21403
rect 14740 21360 14792 21369
rect 15568 21496 15620 21548
rect 19432 21496 19484 21548
rect 20352 21564 20404 21616
rect 20996 21564 21048 21616
rect 21548 21564 21600 21616
rect 21088 21539 21140 21548
rect 21088 21505 21097 21539
rect 21097 21505 21131 21539
rect 21131 21505 21140 21539
rect 21088 21496 21140 21505
rect 22284 21632 22336 21684
rect 15108 21428 15160 21480
rect 16948 21428 17000 21480
rect 18144 21471 18196 21480
rect 18144 21437 18153 21471
rect 18153 21437 18187 21471
rect 18187 21437 18196 21471
rect 18144 21428 18196 21437
rect 19524 21471 19576 21480
rect 19524 21437 19533 21471
rect 19533 21437 19567 21471
rect 19567 21437 19576 21471
rect 19524 21428 19576 21437
rect 19708 21471 19760 21480
rect 19708 21437 19721 21471
rect 19721 21437 19760 21471
rect 19708 21428 19760 21437
rect 20904 21428 20956 21480
rect 21364 21471 21416 21480
rect 21364 21437 21373 21471
rect 21373 21437 21407 21471
rect 21407 21437 21416 21471
rect 21364 21428 21416 21437
rect 21640 21428 21692 21480
rect 21916 21428 21968 21480
rect 15292 21360 15344 21412
rect 16028 21403 16080 21412
rect 16028 21369 16037 21403
rect 16037 21369 16071 21403
rect 16071 21369 16080 21403
rect 16028 21360 16080 21369
rect 15568 21292 15620 21344
rect 15936 21292 15988 21344
rect 17224 21403 17276 21412
rect 17224 21369 17233 21403
rect 17233 21369 17267 21403
rect 17267 21369 17276 21403
rect 17224 21360 17276 21369
rect 17040 21292 17092 21344
rect 17868 21403 17920 21412
rect 17868 21369 17877 21403
rect 17877 21369 17911 21403
rect 17911 21369 17920 21403
rect 17868 21360 17920 21369
rect 19248 21360 19300 21412
rect 18052 21335 18104 21344
rect 18052 21301 18061 21335
rect 18061 21301 18095 21335
rect 18095 21301 18104 21335
rect 18052 21292 18104 21301
rect 18236 21335 18288 21344
rect 18236 21301 18245 21335
rect 18245 21301 18279 21335
rect 18279 21301 18288 21335
rect 18236 21292 18288 21301
rect 19432 21292 19484 21344
rect 20720 21360 20772 21412
rect 21732 21360 21784 21412
rect 20904 21292 20956 21344
rect 21456 21292 21508 21344
rect 4322 21190 4374 21242
rect 4386 21190 4438 21242
rect 4450 21190 4502 21242
rect 4514 21190 4566 21242
rect 4578 21190 4630 21242
rect 4528 21020 4580 21072
rect 4252 20952 4304 21004
rect 7104 21020 7156 21072
rect 9772 21088 9824 21140
rect 10692 21088 10744 21140
rect 5080 20952 5132 21004
rect 7196 20995 7248 21004
rect 7196 20961 7205 20995
rect 7205 20961 7239 20995
rect 7239 20961 7248 20995
rect 7196 20952 7248 20961
rect 7380 20952 7432 21004
rect 8668 21020 8720 21072
rect 7564 20995 7616 21004
rect 7564 20961 7573 20995
rect 7573 20961 7607 20995
rect 7607 20961 7616 20995
rect 7564 20952 7616 20961
rect 8208 20995 8260 21004
rect 8208 20961 8217 20995
rect 8217 20961 8251 20995
rect 8251 20961 8260 20995
rect 8208 20952 8260 20961
rect 8484 20995 8536 21004
rect 8484 20961 8493 20995
rect 8493 20961 8527 20995
rect 8527 20961 8536 20995
rect 8944 20995 8996 21004
rect 8484 20952 8536 20961
rect 8944 20961 8953 20995
rect 8953 20961 8987 20995
rect 8987 20961 8996 20995
rect 8944 20952 8996 20961
rect 9128 20995 9180 21004
rect 9128 20961 9137 20995
rect 9137 20961 9171 20995
rect 9171 20961 9180 20995
rect 9128 20952 9180 20961
rect 9220 20995 9272 21004
rect 9220 20961 9229 20995
rect 9229 20961 9263 20995
rect 9263 20961 9272 20995
rect 9220 20952 9272 20961
rect 9312 20952 9364 21004
rect 10140 21020 10192 21072
rect 14188 21088 14240 21140
rect 15016 21088 15068 21140
rect 15568 21088 15620 21140
rect 17224 21088 17276 21140
rect 10048 20995 10100 21004
rect 10048 20961 10057 20995
rect 10057 20961 10091 20995
rect 10091 20961 10100 20995
rect 10048 20952 10100 20961
rect 12256 20995 12308 21004
rect 12256 20961 12265 20995
rect 12265 20961 12299 20995
rect 12299 20961 12308 20995
rect 12256 20952 12308 20961
rect 6368 20884 6420 20936
rect 14832 21020 14884 21072
rect 12808 20952 12860 21004
rect 13084 20995 13136 21004
rect 13084 20961 13093 20995
rect 13093 20961 13127 20995
rect 13127 20961 13136 20995
rect 13084 20952 13136 20961
rect 14740 20995 14792 21004
rect 14740 20961 14749 20995
rect 14749 20961 14783 20995
rect 14783 20961 14792 20995
rect 14740 20952 14792 20961
rect 10692 20816 10744 20868
rect 14188 20884 14240 20936
rect 15568 20995 15620 21004
rect 15568 20961 15577 20995
rect 15577 20961 15611 20995
rect 15611 20961 15620 20995
rect 15568 20952 15620 20961
rect 16028 21020 16080 21072
rect 17040 21063 17092 21072
rect 17040 21029 17049 21063
rect 17049 21029 17083 21063
rect 17083 21029 17092 21063
rect 17040 21020 17092 21029
rect 15936 20995 15988 21004
rect 15936 20961 15945 20995
rect 15945 20961 15979 20995
rect 15979 20961 15988 20995
rect 15936 20952 15988 20961
rect 16764 20995 16816 21004
rect 16764 20961 16773 20995
rect 16773 20961 16807 20995
rect 16807 20961 16816 20995
rect 16764 20952 16816 20961
rect 18236 20952 18288 21004
rect 19524 20995 19576 21004
rect 19524 20961 19563 20995
rect 19563 20961 19576 20995
rect 19524 20952 19576 20961
rect 19708 20995 19760 21004
rect 19708 20961 19717 20995
rect 19717 20961 19751 20995
rect 19751 20961 19760 20995
rect 19708 20952 19760 20961
rect 20628 20952 20680 21004
rect 21732 20995 21784 21004
rect 21732 20961 21741 20995
rect 21741 20961 21775 20995
rect 21775 20961 21784 20995
rect 21732 20952 21784 20961
rect 16304 20816 16356 20868
rect 18052 20884 18104 20936
rect 17868 20816 17920 20868
rect 20996 20816 21048 20868
rect 21548 20927 21600 20936
rect 21548 20893 21557 20927
rect 21557 20893 21591 20927
rect 21591 20893 21600 20927
rect 21548 20884 21600 20893
rect 22100 20859 22152 20868
rect 9036 20748 9088 20800
rect 9404 20748 9456 20800
rect 11152 20748 11204 20800
rect 12808 20748 12860 20800
rect 16212 20791 16264 20800
rect 16212 20757 16221 20791
rect 16221 20757 16255 20791
rect 16255 20757 16264 20791
rect 16212 20748 16264 20757
rect 17776 20791 17828 20800
rect 17776 20757 17785 20791
rect 17785 20757 17819 20791
rect 17819 20757 17828 20791
rect 17776 20748 17828 20757
rect 19616 20748 19668 20800
rect 21272 20791 21324 20800
rect 21272 20757 21281 20791
rect 21281 20757 21315 20791
rect 21315 20757 21324 20791
rect 21272 20748 21324 20757
rect 22100 20825 22109 20859
rect 22109 20825 22143 20859
rect 22143 20825 22152 20859
rect 22100 20816 22152 20825
rect 21548 20748 21600 20800
rect 3662 20646 3714 20698
rect 3726 20646 3778 20698
rect 3790 20646 3842 20698
rect 3854 20646 3906 20698
rect 3918 20646 3970 20698
rect 4528 20544 4580 20596
rect 5264 20544 5316 20596
rect 10048 20544 10100 20596
rect 10968 20544 11020 20596
rect 4804 20476 4856 20528
rect 4620 20340 4672 20392
rect 4068 20272 4120 20324
rect 4988 20383 5040 20392
rect 4988 20349 4997 20383
rect 4997 20349 5031 20383
rect 5031 20349 5040 20383
rect 4988 20340 5040 20349
rect 5264 20383 5316 20392
rect 5264 20349 5273 20383
rect 5273 20349 5307 20383
rect 5307 20349 5316 20383
rect 5264 20340 5316 20349
rect 6276 20408 6328 20460
rect 5540 20383 5592 20392
rect 5540 20349 5549 20383
rect 5549 20349 5583 20383
rect 5583 20349 5592 20383
rect 5540 20340 5592 20349
rect 7380 20340 7432 20392
rect 9036 20340 9088 20392
rect 9588 20340 9640 20392
rect 15108 20340 15160 20392
rect 16672 20340 16724 20392
rect 19432 20383 19484 20392
rect 19432 20349 19441 20383
rect 19441 20349 19475 20383
rect 19475 20349 19484 20383
rect 19432 20340 19484 20349
rect 19616 20383 19668 20392
rect 19616 20349 19625 20383
rect 19625 20349 19659 20383
rect 19659 20349 19668 20383
rect 19616 20340 19668 20349
rect 20444 20340 20496 20392
rect 21456 20476 21508 20528
rect 20628 20408 20680 20460
rect 20720 20340 20772 20392
rect 4896 20315 4948 20324
rect 4896 20281 4905 20315
rect 4905 20281 4939 20315
rect 4939 20281 4948 20315
rect 4896 20272 4948 20281
rect 14740 20272 14792 20324
rect 20628 20315 20680 20324
rect 20628 20281 20637 20315
rect 20637 20281 20671 20315
rect 20671 20281 20680 20315
rect 20628 20272 20680 20281
rect 20996 20272 21048 20324
rect 6736 20204 6788 20256
rect 19156 20204 19208 20256
rect 20720 20204 20772 20256
rect 21548 20315 21600 20324
rect 21548 20281 21575 20315
rect 21575 20281 21600 20315
rect 21548 20272 21600 20281
rect 4322 20102 4374 20154
rect 4386 20102 4438 20154
rect 4450 20102 4502 20154
rect 4514 20102 4566 20154
rect 4578 20102 4630 20154
rect 2872 19932 2924 19984
rect 2780 19907 2832 19916
rect 2780 19873 2789 19907
rect 2789 19873 2823 19907
rect 2823 19873 2832 19907
rect 2780 19864 2832 19873
rect 3332 19932 3384 19984
rect 4068 19932 4120 19984
rect 5080 20000 5132 20052
rect 21272 20043 21324 20052
rect 21272 20009 21281 20043
rect 21281 20009 21315 20043
rect 21315 20009 21324 20043
rect 21272 20000 21324 20009
rect 4988 19932 5040 19984
rect 3424 19864 3476 19916
rect 4896 19907 4948 19916
rect 4896 19873 4905 19907
rect 4905 19873 4939 19907
rect 4939 19873 4948 19907
rect 4896 19864 4948 19873
rect 8760 19864 8812 19916
rect 9128 19907 9180 19916
rect 9128 19873 9137 19907
rect 9137 19873 9171 19907
rect 9171 19873 9180 19907
rect 9128 19864 9180 19873
rect 9864 19907 9916 19916
rect 9864 19873 9873 19907
rect 9873 19873 9907 19907
rect 9907 19873 9916 19907
rect 9864 19864 9916 19873
rect 9496 19796 9548 19848
rect 4896 19728 4948 19780
rect 11244 19864 11296 19916
rect 18696 19864 18748 19916
rect 19064 19907 19116 19916
rect 19064 19873 19073 19907
rect 19073 19873 19107 19907
rect 19107 19873 19116 19907
rect 19064 19864 19116 19873
rect 19156 19907 19208 19916
rect 19156 19873 19165 19907
rect 19165 19873 19199 19907
rect 19199 19873 19208 19907
rect 19156 19864 19208 19873
rect 19340 19864 19392 19916
rect 20996 19907 21048 19916
rect 20996 19873 21005 19907
rect 21005 19873 21039 19907
rect 21039 19873 21048 19907
rect 20996 19864 21048 19873
rect 21640 19907 21692 19916
rect 21640 19873 21649 19907
rect 21649 19873 21683 19907
rect 21683 19873 21692 19907
rect 21640 19864 21692 19873
rect 11060 19839 11112 19848
rect 11060 19805 11069 19839
rect 11069 19805 11103 19839
rect 11103 19805 11112 19839
rect 11060 19796 11112 19805
rect 21364 19796 21416 19848
rect 3148 19703 3200 19712
rect 3148 19669 3157 19703
rect 3157 19669 3191 19703
rect 3191 19669 3200 19703
rect 3148 19660 3200 19669
rect 3240 19660 3292 19712
rect 6000 19660 6052 19712
rect 7656 19703 7708 19712
rect 7656 19669 7665 19703
rect 7665 19669 7699 19703
rect 7699 19669 7708 19703
rect 7656 19660 7708 19669
rect 11520 19703 11572 19712
rect 11520 19669 11529 19703
rect 11529 19669 11563 19703
rect 11563 19669 11572 19703
rect 11520 19660 11572 19669
rect 19432 19660 19484 19712
rect 19616 19660 19668 19712
rect 20352 19703 20404 19712
rect 20352 19669 20361 19703
rect 20361 19669 20395 19703
rect 20395 19669 20404 19703
rect 20352 19660 20404 19669
rect 20536 19660 20588 19712
rect 3662 19558 3714 19610
rect 3726 19558 3778 19610
rect 3790 19558 3842 19610
rect 3854 19558 3906 19610
rect 3918 19558 3970 19610
rect 2872 19431 2924 19440
rect 2872 19397 2881 19431
rect 2881 19397 2915 19431
rect 2915 19397 2924 19431
rect 2872 19388 2924 19397
rect 3148 19388 3200 19440
rect 3700 19388 3752 19440
rect 5448 19456 5500 19508
rect 2780 19252 2832 19304
rect 3332 19295 3384 19304
rect 3332 19261 3341 19295
rect 3341 19261 3375 19295
rect 3375 19261 3384 19295
rect 3332 19252 3384 19261
rect 4896 19363 4948 19372
rect 4896 19329 4905 19363
rect 4905 19329 4939 19363
rect 4939 19329 4948 19363
rect 4896 19320 4948 19329
rect 7196 19388 7248 19440
rect 7656 19388 7708 19440
rect 6736 19363 6788 19372
rect 6736 19329 6745 19363
rect 6745 19329 6779 19363
rect 6779 19329 6788 19363
rect 6736 19320 6788 19329
rect 3608 19295 3660 19304
rect 3608 19261 3617 19295
rect 3617 19261 3651 19295
rect 3651 19261 3660 19295
rect 3608 19252 3660 19261
rect 3516 19184 3568 19236
rect 4988 19295 5040 19304
rect 4988 19261 4997 19295
rect 4997 19261 5031 19295
rect 5031 19261 5040 19295
rect 4988 19252 5040 19261
rect 6000 19295 6052 19304
rect 6000 19261 6009 19295
rect 6009 19261 6043 19295
rect 6043 19261 6052 19295
rect 6000 19252 6052 19261
rect 7380 19320 7432 19372
rect 11520 19320 11572 19372
rect 12164 19320 12216 19372
rect 8392 19252 8444 19304
rect 8760 19252 8812 19304
rect 4252 19159 4304 19168
rect 4252 19125 4261 19159
rect 4261 19125 4295 19159
rect 4295 19125 4304 19159
rect 4252 19116 4304 19125
rect 6276 19159 6328 19168
rect 6276 19125 6285 19159
rect 6285 19125 6319 19159
rect 6319 19125 6328 19159
rect 6276 19116 6328 19125
rect 9496 19184 9548 19236
rect 9772 19184 9824 19236
rect 10692 19295 10744 19304
rect 10692 19261 10701 19295
rect 10701 19261 10735 19295
rect 10735 19261 10744 19295
rect 10692 19252 10744 19261
rect 10968 19252 11020 19304
rect 12992 19295 13044 19304
rect 12992 19261 13001 19295
rect 13001 19261 13035 19295
rect 13035 19261 13044 19295
rect 12992 19252 13044 19261
rect 13176 19320 13228 19372
rect 17592 19456 17644 19508
rect 13268 19252 13320 19304
rect 16212 19252 16264 19304
rect 17776 19320 17828 19372
rect 10600 19184 10652 19236
rect 15200 19184 15252 19236
rect 7104 19116 7156 19168
rect 7564 19159 7616 19168
rect 7564 19125 7573 19159
rect 7573 19125 7607 19159
rect 7607 19125 7616 19159
rect 7564 19116 7616 19125
rect 16396 19159 16448 19168
rect 16396 19125 16405 19159
rect 16405 19125 16439 19159
rect 16439 19125 16448 19159
rect 17132 19295 17184 19304
rect 17132 19261 17141 19295
rect 17141 19261 17175 19295
rect 17175 19261 17184 19295
rect 17132 19252 17184 19261
rect 17316 19227 17368 19236
rect 17316 19193 17325 19227
rect 17325 19193 17359 19227
rect 17359 19193 17368 19227
rect 17316 19184 17368 19193
rect 17776 19184 17828 19236
rect 17960 19295 18012 19304
rect 17960 19261 17969 19295
rect 17969 19261 18003 19295
rect 18003 19261 18012 19295
rect 17960 19252 18012 19261
rect 20352 19388 20404 19440
rect 19432 19363 19484 19372
rect 19432 19329 19441 19363
rect 19441 19329 19475 19363
rect 19475 19329 19484 19363
rect 19432 19320 19484 19329
rect 18696 19295 18748 19304
rect 18696 19261 18705 19295
rect 18705 19261 18739 19295
rect 18739 19261 18748 19295
rect 18696 19252 18748 19261
rect 19156 19252 19208 19304
rect 18420 19184 18472 19236
rect 19616 19295 19668 19304
rect 19616 19261 19625 19295
rect 19625 19261 19659 19295
rect 19659 19261 19668 19295
rect 19616 19252 19668 19261
rect 19708 19295 19760 19304
rect 19708 19261 19717 19295
rect 19717 19261 19751 19295
rect 19751 19261 19760 19295
rect 19708 19252 19760 19261
rect 20352 19295 20404 19304
rect 20352 19261 20361 19295
rect 20361 19261 20395 19295
rect 20395 19261 20404 19295
rect 20352 19252 20404 19261
rect 20536 19295 20588 19304
rect 20536 19261 20545 19295
rect 20545 19261 20579 19295
rect 20579 19261 20588 19295
rect 20536 19252 20588 19261
rect 20812 19252 20864 19304
rect 21088 19295 21140 19304
rect 21088 19261 21097 19295
rect 21097 19261 21131 19295
rect 21131 19261 21140 19295
rect 21088 19252 21140 19261
rect 21364 19252 21416 19304
rect 21456 19295 21508 19304
rect 21456 19261 21468 19295
rect 21468 19261 21502 19295
rect 21502 19261 21508 19295
rect 21456 19252 21508 19261
rect 22284 19295 22336 19304
rect 22284 19261 22293 19295
rect 22293 19261 22327 19295
rect 22327 19261 22336 19295
rect 22284 19252 22336 19261
rect 22376 19295 22428 19304
rect 22376 19261 22385 19295
rect 22385 19261 22419 19295
rect 22419 19261 22428 19295
rect 22376 19252 22428 19261
rect 22560 19295 22612 19304
rect 22560 19261 22569 19295
rect 22569 19261 22603 19295
rect 22603 19261 22612 19295
rect 22560 19252 22612 19261
rect 23020 19295 23072 19304
rect 23020 19261 23029 19295
rect 23029 19261 23063 19295
rect 23063 19261 23072 19295
rect 23020 19252 23072 19261
rect 16396 19116 16448 19125
rect 18052 19116 18104 19168
rect 18144 19116 18196 19168
rect 19064 19116 19116 19168
rect 20444 19184 20496 19236
rect 21180 19184 21232 19236
rect 19248 19159 19300 19168
rect 19248 19125 19257 19159
rect 19257 19125 19291 19159
rect 19291 19125 19300 19159
rect 19248 19116 19300 19125
rect 21364 19116 21416 19168
rect 21640 19159 21692 19168
rect 21640 19125 21649 19159
rect 21649 19125 21683 19159
rect 21683 19125 21692 19159
rect 21640 19116 21692 19125
rect 4322 19014 4374 19066
rect 4386 19014 4438 19066
rect 4450 19014 4502 19066
rect 4514 19014 4566 19066
rect 4578 19014 4630 19066
rect 3608 18912 3660 18964
rect 5264 18912 5316 18964
rect 2780 18887 2832 18896
rect 2780 18853 2789 18887
rect 2789 18853 2823 18887
rect 2823 18853 2832 18887
rect 2780 18844 2832 18853
rect 5540 18844 5592 18896
rect 3700 18819 3752 18828
rect 3700 18785 3709 18819
rect 3709 18785 3743 18819
rect 3743 18785 3752 18819
rect 3700 18776 3752 18785
rect 4160 18819 4212 18828
rect 4160 18785 4169 18819
rect 4169 18785 4203 18819
rect 4203 18785 4212 18819
rect 4160 18776 4212 18785
rect 4988 18819 5040 18828
rect 4988 18785 4997 18819
rect 4997 18785 5031 18819
rect 5031 18785 5040 18819
rect 4988 18776 5040 18785
rect 6276 18844 6328 18896
rect 5080 18751 5132 18760
rect 5080 18717 5089 18751
rect 5089 18717 5123 18751
rect 5123 18717 5132 18751
rect 5080 18708 5132 18717
rect 5448 18708 5500 18760
rect 6644 18819 6696 18828
rect 6644 18785 6653 18819
rect 6653 18785 6687 18819
rect 6687 18785 6696 18819
rect 6644 18776 6696 18785
rect 7288 18776 7340 18828
rect 9036 18844 9088 18896
rect 10692 18844 10744 18896
rect 10968 18844 11020 18896
rect 12256 18912 12308 18964
rect 15292 18912 15344 18964
rect 3240 18640 3292 18692
rect 4896 18640 4948 18692
rect 7380 18708 7432 18760
rect 6828 18640 6880 18692
rect 6920 18640 6972 18692
rect 7564 18751 7616 18760
rect 7564 18717 7573 18751
rect 7573 18717 7607 18751
rect 7607 18717 7616 18751
rect 8760 18776 8812 18828
rect 9588 18819 9640 18828
rect 9588 18785 9597 18819
rect 9597 18785 9631 18819
rect 9631 18785 9640 18819
rect 9588 18776 9640 18785
rect 10416 18819 10468 18828
rect 10416 18785 10425 18819
rect 10425 18785 10459 18819
rect 10459 18785 10468 18819
rect 10416 18776 10468 18785
rect 10600 18819 10652 18828
rect 10600 18785 10609 18819
rect 10609 18785 10643 18819
rect 10643 18785 10652 18819
rect 10600 18776 10652 18785
rect 11060 18776 11112 18828
rect 12164 18819 12216 18828
rect 12164 18785 12173 18819
rect 12173 18785 12207 18819
rect 12207 18785 12216 18819
rect 12164 18776 12216 18785
rect 12716 18819 12768 18828
rect 12716 18785 12725 18819
rect 12725 18785 12759 18819
rect 12759 18785 12768 18819
rect 12716 18776 12768 18785
rect 12992 18819 13044 18828
rect 12992 18785 13001 18819
rect 13001 18785 13035 18819
rect 13035 18785 13044 18819
rect 12992 18776 13044 18785
rect 13360 18776 13412 18828
rect 15752 18776 15804 18828
rect 17316 18912 17368 18964
rect 17960 18912 18012 18964
rect 18420 18955 18472 18964
rect 18420 18921 18429 18955
rect 18429 18921 18463 18955
rect 18463 18921 18472 18955
rect 18420 18912 18472 18921
rect 20352 18912 20404 18964
rect 21456 18912 21508 18964
rect 17776 18844 17828 18896
rect 19248 18844 19300 18896
rect 21640 18844 21692 18896
rect 17224 18819 17276 18828
rect 7564 18708 7616 18717
rect 8484 18708 8536 18760
rect 11244 18751 11296 18760
rect 11244 18717 11253 18751
rect 11253 18717 11287 18751
rect 11287 18717 11296 18751
rect 11244 18708 11296 18717
rect 12532 18708 12584 18760
rect 13268 18708 13320 18760
rect 14556 18751 14608 18760
rect 14556 18717 14565 18751
rect 14565 18717 14599 18751
rect 14599 18717 14608 18751
rect 14556 18708 14608 18717
rect 16396 18751 16448 18760
rect 16396 18717 16405 18751
rect 16405 18717 16439 18751
rect 16439 18717 16448 18751
rect 16396 18708 16448 18717
rect 17224 18785 17233 18819
rect 17233 18785 17267 18819
rect 17267 18785 17276 18819
rect 17224 18776 17276 18785
rect 17408 18819 17460 18828
rect 17408 18785 17417 18819
rect 17417 18785 17451 18819
rect 17451 18785 17460 18819
rect 17408 18776 17460 18785
rect 17592 18819 17644 18828
rect 17592 18785 17601 18819
rect 17601 18785 17635 18819
rect 17635 18785 17644 18819
rect 17592 18776 17644 18785
rect 18052 18819 18104 18828
rect 18052 18785 18061 18819
rect 18061 18785 18095 18819
rect 18095 18785 18104 18819
rect 18052 18776 18104 18785
rect 17132 18708 17184 18760
rect 3516 18572 3568 18624
rect 4068 18572 4120 18624
rect 9496 18640 9548 18692
rect 13912 18640 13964 18692
rect 19616 18776 19668 18828
rect 21272 18776 21324 18828
rect 18880 18751 18932 18760
rect 18880 18717 18889 18751
rect 18889 18717 18923 18751
rect 18923 18717 18932 18751
rect 18880 18708 18932 18717
rect 20904 18708 20956 18760
rect 22652 18751 22704 18760
rect 22652 18717 22661 18751
rect 22661 18717 22695 18751
rect 22695 18717 22704 18751
rect 22652 18708 22704 18717
rect 8208 18615 8260 18624
rect 8208 18581 8217 18615
rect 8217 18581 8251 18615
rect 8251 18581 8260 18615
rect 8208 18572 8260 18581
rect 8300 18615 8352 18624
rect 8300 18581 8309 18615
rect 8309 18581 8343 18615
rect 8343 18581 8352 18615
rect 8300 18572 8352 18581
rect 10048 18572 10100 18624
rect 12624 18572 12676 18624
rect 12900 18615 12952 18624
rect 12900 18581 12909 18615
rect 12909 18581 12943 18615
rect 12943 18581 12952 18615
rect 12900 18572 12952 18581
rect 15016 18615 15068 18624
rect 15016 18581 15025 18615
rect 15025 18581 15059 18615
rect 15059 18581 15068 18615
rect 15016 18572 15068 18581
rect 17776 18572 17828 18624
rect 18420 18572 18472 18624
rect 20076 18572 20128 18624
rect 21088 18572 21140 18624
rect 21640 18572 21692 18624
rect 22284 18572 22336 18624
rect 3662 18470 3714 18522
rect 3726 18470 3778 18522
rect 3790 18470 3842 18522
rect 3854 18470 3906 18522
rect 3918 18470 3970 18522
rect 6276 18368 6328 18420
rect 12624 18411 12676 18420
rect 12624 18377 12633 18411
rect 12633 18377 12667 18411
rect 12667 18377 12676 18411
rect 12624 18368 12676 18377
rect 9588 18300 9640 18352
rect 10048 18300 10100 18352
rect 3332 18232 3384 18284
rect 4252 18232 4304 18284
rect 7380 18232 7432 18284
rect 4344 18164 4396 18216
rect 4896 18164 4948 18216
rect 5264 18207 5316 18216
rect 5264 18173 5273 18207
rect 5273 18173 5307 18207
rect 5307 18173 5316 18207
rect 5264 18164 5316 18173
rect 7288 18207 7340 18216
rect 7288 18173 7297 18207
rect 7297 18173 7331 18207
rect 7331 18173 7340 18207
rect 7288 18164 7340 18173
rect 7472 18207 7524 18216
rect 7472 18173 7481 18207
rect 7481 18173 7515 18207
rect 7515 18173 7524 18207
rect 7472 18164 7524 18173
rect 9956 18232 10008 18284
rect 8392 18164 8444 18216
rect 8760 18207 8812 18216
rect 8760 18173 8769 18207
rect 8769 18173 8803 18207
rect 8803 18173 8812 18207
rect 8760 18164 8812 18173
rect 5080 18139 5132 18148
rect 5080 18105 5089 18139
rect 5089 18105 5123 18139
rect 5123 18105 5132 18139
rect 5080 18096 5132 18105
rect 9036 18096 9088 18148
rect 10048 18207 10100 18216
rect 10048 18173 10057 18207
rect 10057 18173 10091 18207
rect 10091 18173 10100 18207
rect 10048 18164 10100 18173
rect 10416 18164 10468 18216
rect 10692 18164 10744 18216
rect 11152 18207 11204 18216
rect 11152 18173 11161 18207
rect 11161 18173 11195 18207
rect 11195 18173 11204 18207
rect 11152 18164 11204 18173
rect 12440 18300 12492 18352
rect 19708 18411 19760 18420
rect 19708 18377 19717 18411
rect 19717 18377 19751 18411
rect 19751 18377 19760 18411
rect 19708 18368 19760 18377
rect 20996 18411 21048 18420
rect 20996 18377 21005 18411
rect 21005 18377 21039 18411
rect 21039 18377 21048 18411
rect 20996 18368 21048 18377
rect 21180 18368 21232 18420
rect 22284 18368 22336 18420
rect 13084 18300 13136 18352
rect 12716 18232 12768 18284
rect 12532 18207 12584 18216
rect 12532 18173 12541 18207
rect 12541 18173 12575 18207
rect 12575 18173 12584 18207
rect 12532 18164 12584 18173
rect 13268 18232 13320 18284
rect 14924 18300 14976 18352
rect 15292 18300 15344 18352
rect 15016 18232 15068 18284
rect 11060 18096 11112 18148
rect 12256 18096 12308 18148
rect 7380 18071 7432 18080
rect 7380 18037 7389 18071
rect 7389 18037 7423 18071
rect 7423 18037 7432 18071
rect 7380 18028 7432 18037
rect 7748 18071 7800 18080
rect 7748 18037 7757 18071
rect 7757 18037 7791 18071
rect 7791 18037 7800 18071
rect 7748 18028 7800 18037
rect 12164 18028 12216 18080
rect 13452 18096 13504 18148
rect 15292 18207 15344 18216
rect 15292 18173 15301 18207
rect 15301 18173 15335 18207
rect 15335 18173 15344 18207
rect 15292 18164 15344 18173
rect 15752 18207 15804 18216
rect 15752 18173 15761 18207
rect 15761 18173 15795 18207
rect 15795 18173 15804 18207
rect 15752 18164 15804 18173
rect 17224 18275 17276 18284
rect 17224 18241 17233 18275
rect 17233 18241 17267 18275
rect 17267 18241 17276 18275
rect 17224 18232 17276 18241
rect 20812 18232 20864 18284
rect 17408 18207 17460 18216
rect 14556 18096 14608 18148
rect 17408 18173 17417 18207
rect 17417 18173 17451 18207
rect 17451 18173 17460 18207
rect 17408 18164 17460 18173
rect 19892 18207 19944 18216
rect 19892 18173 19901 18207
rect 19901 18173 19935 18207
rect 19935 18173 19944 18207
rect 19892 18164 19944 18173
rect 20076 18207 20128 18216
rect 20076 18173 20085 18207
rect 20085 18173 20119 18207
rect 20119 18173 20128 18207
rect 20076 18164 20128 18173
rect 21364 18232 21416 18284
rect 21640 18207 21692 18216
rect 21640 18173 21649 18207
rect 21649 18173 21683 18207
rect 21683 18173 21692 18207
rect 21640 18164 21692 18173
rect 18880 18096 18932 18148
rect 13912 18028 13964 18080
rect 14004 18071 14056 18080
rect 14004 18037 14013 18071
rect 14013 18037 14047 18071
rect 14047 18037 14056 18071
rect 14004 18028 14056 18037
rect 15660 18071 15712 18080
rect 15660 18037 15669 18071
rect 15669 18037 15703 18071
rect 15703 18037 15712 18071
rect 15660 18028 15712 18037
rect 17684 18028 17736 18080
rect 4322 17926 4374 17978
rect 4386 17926 4438 17978
rect 4450 17926 4502 17978
rect 4514 17926 4566 17978
rect 4578 17926 4630 17978
rect 5080 17824 5132 17876
rect 11152 17824 11204 17876
rect 15292 17824 15344 17876
rect 2780 17756 2832 17808
rect 3424 17756 3476 17808
rect 3332 17688 3384 17740
rect 9496 17756 9548 17808
rect 3148 17620 3200 17672
rect 9588 17731 9640 17740
rect 9588 17697 9597 17731
rect 9597 17697 9631 17731
rect 9631 17697 9640 17731
rect 9588 17688 9640 17697
rect 12440 17688 12492 17740
rect 13452 17756 13504 17808
rect 13912 17756 13964 17808
rect 13176 17731 13228 17740
rect 13176 17697 13185 17731
rect 13185 17697 13219 17731
rect 13219 17697 13228 17731
rect 13176 17688 13228 17697
rect 14004 17688 14056 17740
rect 22100 17756 22152 17808
rect 22836 17756 22888 17808
rect 17684 17731 17736 17740
rect 17684 17697 17693 17731
rect 17693 17697 17727 17731
rect 17727 17697 17736 17731
rect 17684 17688 17736 17697
rect 17776 17688 17828 17740
rect 21640 17731 21692 17740
rect 21640 17697 21649 17731
rect 21649 17697 21683 17731
rect 21683 17697 21692 17731
rect 21640 17688 21692 17697
rect 22008 17688 22060 17740
rect 9496 17663 9548 17672
rect 9496 17629 9505 17663
rect 9505 17629 9539 17663
rect 9539 17629 9548 17663
rect 9496 17620 9548 17629
rect 9956 17663 10008 17672
rect 9956 17629 9965 17663
rect 9965 17629 9999 17663
rect 9999 17629 10008 17663
rect 9956 17620 10008 17629
rect 13912 17620 13964 17672
rect 12900 17484 12952 17536
rect 14004 17484 14056 17536
rect 14280 17527 14332 17536
rect 14280 17493 14289 17527
rect 14289 17493 14323 17527
rect 14323 17493 14332 17527
rect 14280 17484 14332 17493
rect 17868 17484 17920 17536
rect 21732 17484 21784 17536
rect 3662 17382 3714 17434
rect 3726 17382 3778 17434
rect 3790 17382 3842 17434
rect 3854 17382 3906 17434
rect 3918 17382 3970 17434
rect 3516 17280 3568 17332
rect 9588 17280 9640 17332
rect 9680 17280 9732 17332
rect 14556 17280 14608 17332
rect 18420 17280 18472 17332
rect 7012 17144 7064 17196
rect 8116 17144 8168 17196
rect 13544 17144 13596 17196
rect 14280 17212 14332 17264
rect 14096 17187 14148 17196
rect 14096 17153 14105 17187
rect 14105 17153 14139 17187
rect 14139 17153 14148 17187
rect 14096 17144 14148 17153
rect 5448 17076 5500 17128
rect 6092 17119 6144 17128
rect 6092 17085 6101 17119
rect 6101 17085 6135 17119
rect 6135 17085 6144 17119
rect 6092 17076 6144 17085
rect 8852 17076 8904 17128
rect 13176 17076 13228 17128
rect 13728 17119 13780 17128
rect 13728 17085 13737 17119
rect 13737 17085 13771 17119
rect 13771 17085 13780 17119
rect 13728 17076 13780 17085
rect 3332 17008 3384 17060
rect 3608 17008 3660 17060
rect 13636 17008 13688 17060
rect 16764 17212 16816 17264
rect 15660 17187 15712 17196
rect 15660 17153 15669 17187
rect 15669 17153 15703 17187
rect 15703 17153 15712 17187
rect 15660 17144 15712 17153
rect 17776 17144 17828 17196
rect 17868 17119 17920 17128
rect 17868 17085 17877 17119
rect 17877 17085 17911 17119
rect 17911 17085 17920 17119
rect 17868 17076 17920 17085
rect 18420 17187 18472 17196
rect 18420 17153 18429 17187
rect 18429 17153 18463 17187
rect 18463 17153 18472 17187
rect 18420 17144 18472 17153
rect 18972 17119 19024 17128
rect 18972 17085 18981 17119
rect 18981 17085 19015 17119
rect 19015 17085 19024 17119
rect 18972 17076 19024 17085
rect 19064 17076 19116 17128
rect 19616 17144 19668 17196
rect 20720 17280 20772 17332
rect 22836 17323 22888 17332
rect 22836 17289 22845 17323
rect 22845 17289 22879 17323
rect 22879 17289 22888 17323
rect 22836 17280 22888 17289
rect 18328 17008 18380 17060
rect 18788 17008 18840 17060
rect 3424 16940 3476 16992
rect 4068 16983 4120 16992
rect 4068 16949 4077 16983
rect 4077 16949 4111 16983
rect 4111 16949 4120 16983
rect 4068 16940 4120 16949
rect 7472 16940 7524 16992
rect 11520 16940 11572 16992
rect 15108 16940 15160 16992
rect 16028 16983 16080 16992
rect 16028 16949 16037 16983
rect 16037 16949 16071 16983
rect 16071 16949 16080 16983
rect 16028 16940 16080 16949
rect 17960 16983 18012 16992
rect 17960 16949 17969 16983
rect 17969 16949 18003 16983
rect 18003 16949 18012 16983
rect 17960 16940 18012 16949
rect 18696 16983 18748 16992
rect 18696 16949 18705 16983
rect 18705 16949 18739 16983
rect 18739 16949 18748 16983
rect 18696 16940 18748 16949
rect 20444 17119 20496 17128
rect 20444 17085 20453 17119
rect 20453 17085 20487 17119
rect 20487 17085 20496 17119
rect 20444 17076 20496 17085
rect 22376 17076 22428 17128
rect 22836 17076 22888 17128
rect 22192 17051 22244 17060
rect 22192 17017 22201 17051
rect 22201 17017 22235 17051
rect 22235 17017 22244 17051
rect 22192 17008 22244 17017
rect 21456 16940 21508 16992
rect 22744 16940 22796 16992
rect 4322 16838 4374 16890
rect 4386 16838 4438 16890
rect 4450 16838 4502 16890
rect 4514 16838 4566 16890
rect 4578 16838 4630 16890
rect 4160 16736 4212 16788
rect 5448 16736 5500 16788
rect 9680 16736 9732 16788
rect 11520 16779 11572 16788
rect 11520 16745 11529 16779
rect 11529 16745 11563 16779
rect 11563 16745 11572 16779
rect 11520 16736 11572 16745
rect 12348 16736 12400 16788
rect 15384 16736 15436 16788
rect 2872 16643 2924 16652
rect 2872 16609 2881 16643
rect 2881 16609 2915 16643
rect 2915 16609 2924 16643
rect 2872 16600 2924 16609
rect 3148 16643 3200 16652
rect 3148 16609 3157 16643
rect 3157 16609 3191 16643
rect 3191 16609 3200 16643
rect 3148 16600 3200 16609
rect 3056 16532 3108 16584
rect 3516 16643 3568 16652
rect 3516 16609 3525 16643
rect 3525 16609 3559 16643
rect 3559 16609 3568 16643
rect 3516 16600 3568 16609
rect 3884 16600 3936 16652
rect 4068 16600 4120 16652
rect 7012 16668 7064 16720
rect 7748 16668 7800 16720
rect 8116 16668 8168 16720
rect 8300 16668 8352 16720
rect 4620 16532 4672 16584
rect 5264 16600 5316 16652
rect 6276 16643 6328 16652
rect 6276 16609 6285 16643
rect 6285 16609 6319 16643
rect 6319 16609 6328 16643
rect 6276 16600 6328 16609
rect 7104 16600 7156 16652
rect 7472 16643 7524 16652
rect 7472 16609 7481 16643
rect 7481 16609 7515 16643
rect 7515 16609 7524 16643
rect 7472 16600 7524 16609
rect 11060 16668 11112 16720
rect 13636 16668 13688 16720
rect 14004 16711 14056 16720
rect 14004 16677 14013 16711
rect 14013 16677 14047 16711
rect 14047 16677 14056 16711
rect 14004 16668 14056 16677
rect 6460 16575 6512 16584
rect 6460 16541 6469 16575
rect 6469 16541 6503 16575
rect 6503 16541 6512 16575
rect 6460 16532 6512 16541
rect 3516 16464 3568 16516
rect 9680 16532 9732 16584
rect 10968 16575 11020 16584
rect 10968 16541 10977 16575
rect 10977 16541 11011 16575
rect 11011 16541 11020 16575
rect 10968 16532 11020 16541
rect 7748 16464 7800 16516
rect 8852 16464 8904 16516
rect 12164 16600 12216 16652
rect 13728 16643 13780 16652
rect 13728 16609 13737 16643
rect 13737 16609 13771 16643
rect 13771 16609 13780 16643
rect 13728 16600 13780 16609
rect 13912 16600 13964 16652
rect 15200 16668 15252 16720
rect 12348 16575 12400 16584
rect 12348 16541 12357 16575
rect 12357 16541 12391 16575
rect 12391 16541 12400 16575
rect 12348 16532 12400 16541
rect 15108 16643 15160 16652
rect 15108 16609 15117 16643
rect 15117 16609 15151 16643
rect 15151 16609 15160 16643
rect 15108 16600 15160 16609
rect 15660 16600 15712 16652
rect 16856 16736 16908 16788
rect 18144 16779 18196 16788
rect 18144 16745 18153 16779
rect 18153 16745 18187 16779
rect 18187 16745 18196 16779
rect 18144 16736 18196 16745
rect 18420 16736 18472 16788
rect 18972 16736 19024 16788
rect 19156 16736 19208 16788
rect 22836 16779 22888 16788
rect 22836 16745 22845 16779
rect 22845 16745 22879 16779
rect 22879 16745 22888 16779
rect 22836 16736 22888 16745
rect 16028 16668 16080 16720
rect 15844 16532 15896 16584
rect 17132 16643 17184 16652
rect 17132 16609 17141 16643
rect 17141 16609 17175 16643
rect 17175 16609 17184 16643
rect 17132 16600 17184 16609
rect 17316 16643 17368 16652
rect 17316 16609 17325 16643
rect 17325 16609 17359 16643
rect 17359 16609 17368 16643
rect 17316 16600 17368 16609
rect 16948 16532 17000 16584
rect 17868 16600 17920 16652
rect 18328 16600 18380 16652
rect 18880 16668 18932 16720
rect 20444 16668 20496 16720
rect 19248 16600 19300 16652
rect 21180 16600 21232 16652
rect 22652 16668 22704 16720
rect 21732 16643 21784 16652
rect 21732 16609 21766 16643
rect 21766 16609 21784 16643
rect 21732 16600 21784 16609
rect 18236 16464 18288 16516
rect 8208 16396 8260 16448
rect 8576 16439 8628 16448
rect 8576 16405 8585 16439
rect 8585 16405 8619 16439
rect 8619 16405 8628 16439
rect 8576 16396 8628 16405
rect 16488 16396 16540 16448
rect 3662 16294 3714 16346
rect 3726 16294 3778 16346
rect 3790 16294 3842 16346
rect 3854 16294 3906 16346
rect 3918 16294 3970 16346
rect 3148 16124 3200 16176
rect 3424 16056 3476 16108
rect 3976 16056 4028 16108
rect 4160 16056 4212 16108
rect 6092 16056 6144 16108
rect 7104 16099 7156 16108
rect 7104 16065 7113 16099
rect 7113 16065 7147 16099
rect 7147 16065 7156 16099
rect 7104 16056 7156 16065
rect 7748 16099 7800 16108
rect 7748 16065 7757 16099
rect 7757 16065 7791 16099
rect 7791 16065 7800 16099
rect 7748 16056 7800 16065
rect 3516 15988 3568 16040
rect 4620 16031 4672 16040
rect 4620 15997 4629 16031
rect 4629 15997 4663 16031
rect 4663 15997 4672 16031
rect 4620 15988 4672 15997
rect 5448 15988 5500 16040
rect 6276 16031 6328 16040
rect 6276 15997 6285 16031
rect 6285 15997 6319 16031
rect 6319 15997 6328 16031
rect 6276 15988 6328 15997
rect 6460 16031 6512 16040
rect 6460 15997 6469 16031
rect 6469 15997 6503 16031
rect 6503 15997 6512 16031
rect 6460 15988 6512 15997
rect 7196 16031 7248 16040
rect 7196 15997 7205 16031
rect 7205 15997 7239 16031
rect 7239 15997 7248 16031
rect 7196 15988 7248 15997
rect 9036 16192 9088 16244
rect 9680 16235 9732 16244
rect 9680 16201 9689 16235
rect 9689 16201 9723 16235
rect 9723 16201 9732 16235
rect 9680 16192 9732 16201
rect 10968 16192 11020 16244
rect 13544 16235 13596 16244
rect 13544 16201 13553 16235
rect 13553 16201 13587 16235
rect 13587 16201 13596 16235
rect 13544 16192 13596 16201
rect 15844 16235 15896 16244
rect 15844 16201 15853 16235
rect 15853 16201 15887 16235
rect 15887 16201 15896 16235
rect 15844 16192 15896 16201
rect 15936 16192 15988 16244
rect 16856 16235 16908 16244
rect 16856 16201 16865 16235
rect 16865 16201 16899 16235
rect 16899 16201 16908 16235
rect 16856 16192 16908 16201
rect 8300 16124 8352 16176
rect 12624 16124 12676 16176
rect 17316 16192 17368 16244
rect 17960 16192 18012 16244
rect 19248 16235 19300 16244
rect 19248 16201 19257 16235
rect 19257 16201 19291 16235
rect 19291 16201 19300 16235
rect 19248 16192 19300 16201
rect 21640 16192 21692 16244
rect 22008 16235 22060 16244
rect 22008 16201 22017 16235
rect 22017 16201 22051 16235
rect 22051 16201 22060 16235
rect 22008 16192 22060 16201
rect 18972 16124 19024 16176
rect 8024 16056 8076 16108
rect 8668 15988 8720 16040
rect 8852 16031 8904 16040
rect 8852 15997 8861 16031
rect 8861 15997 8895 16031
rect 8895 15997 8904 16031
rect 8852 15988 8904 15997
rect 9036 16031 9088 16040
rect 9036 15997 9045 16031
rect 9045 15997 9079 16031
rect 9079 15997 9088 16031
rect 9036 15988 9088 15997
rect 14004 16056 14056 16108
rect 16028 16056 16080 16108
rect 19892 16124 19944 16176
rect 22284 16124 22336 16176
rect 2872 15963 2924 15972
rect 2872 15929 2881 15963
rect 2881 15929 2915 15963
rect 2915 15929 2924 15963
rect 2872 15920 2924 15929
rect 2964 15920 3016 15972
rect 3608 15920 3660 15972
rect 3700 15920 3752 15972
rect 10968 15988 11020 16040
rect 12808 15988 12860 16040
rect 13268 15988 13320 16040
rect 13452 15988 13504 16040
rect 13728 16031 13780 16040
rect 13728 15997 13737 16031
rect 13737 15997 13771 16031
rect 13771 15997 13780 16031
rect 13728 15988 13780 15997
rect 13912 16031 13964 16040
rect 13912 15997 13921 16031
rect 13921 15997 13955 16031
rect 13955 15997 13964 16031
rect 13912 15988 13964 15997
rect 15384 15988 15436 16040
rect 3056 15895 3108 15904
rect 3056 15861 3065 15895
rect 3065 15861 3099 15895
rect 3099 15861 3108 15895
rect 3056 15852 3108 15861
rect 3792 15852 3844 15904
rect 6368 15895 6420 15904
rect 6368 15861 6377 15895
rect 6377 15861 6411 15895
rect 6411 15861 6420 15895
rect 6368 15852 6420 15861
rect 11060 15920 11112 15972
rect 11612 15920 11664 15972
rect 16488 16031 16540 16040
rect 16488 15997 16497 16031
rect 16497 15997 16531 16031
rect 16531 15997 16540 16031
rect 16488 15988 16540 15997
rect 16764 16031 16816 16040
rect 16764 15997 16773 16031
rect 16773 15997 16807 16031
rect 16807 15997 16816 16031
rect 16764 15988 16816 15997
rect 16948 15988 17000 16040
rect 17132 16031 17184 16040
rect 17132 15997 17141 16031
rect 17141 15997 17175 16031
rect 17175 15997 17184 16031
rect 17132 15988 17184 15997
rect 17960 16031 18012 16040
rect 17960 15997 17969 16031
rect 17969 15997 18003 16031
rect 18003 15997 18012 16031
rect 17960 15988 18012 15997
rect 18420 16031 18472 16040
rect 18420 15997 18429 16031
rect 18429 15997 18463 16031
rect 18463 15997 18472 16031
rect 18420 15988 18472 15997
rect 18696 16031 18748 16040
rect 18696 15997 18705 16031
rect 18705 15997 18739 16031
rect 18739 15997 18748 16031
rect 18696 15988 18748 15997
rect 18788 15988 18840 16040
rect 19524 15988 19576 16040
rect 21456 16031 21508 16040
rect 21456 15997 21465 16031
rect 21465 15997 21499 16031
rect 21499 15997 21508 16031
rect 21456 15988 21508 15997
rect 21548 16031 21600 16040
rect 21548 15997 21557 16031
rect 21557 15997 21591 16031
rect 21591 15997 21600 16031
rect 21548 15988 21600 15997
rect 16580 15963 16632 15972
rect 8392 15895 8444 15904
rect 8392 15861 8401 15895
rect 8401 15861 8435 15895
rect 8435 15861 8444 15895
rect 8392 15852 8444 15861
rect 13176 15852 13228 15904
rect 13452 15852 13504 15904
rect 13728 15852 13780 15904
rect 16580 15929 16589 15963
rect 16589 15929 16623 15963
rect 16623 15929 16632 15963
rect 16580 15920 16632 15929
rect 19156 15920 19208 15972
rect 22192 16056 22244 16108
rect 22100 16031 22152 16040
rect 22100 15997 22109 16031
rect 22109 15997 22143 16031
rect 22143 15997 22152 16031
rect 22100 15988 22152 15997
rect 18328 15852 18380 15904
rect 18512 15852 18564 15904
rect 21732 15895 21784 15904
rect 21732 15861 21741 15895
rect 21741 15861 21775 15895
rect 21775 15861 21784 15895
rect 21732 15852 21784 15861
rect 4322 15750 4374 15802
rect 4386 15750 4438 15802
rect 4450 15750 4502 15802
rect 4514 15750 4566 15802
rect 4578 15750 4630 15802
rect 3056 15648 3108 15700
rect 3700 15623 3752 15632
rect 3700 15589 3717 15623
rect 3717 15589 3752 15623
rect 3700 15580 3752 15589
rect 3792 15623 3844 15632
rect 3792 15589 3801 15623
rect 3801 15589 3835 15623
rect 3835 15589 3844 15623
rect 3792 15580 3844 15589
rect 8024 15691 8076 15700
rect 8024 15657 8033 15691
rect 8033 15657 8067 15691
rect 8067 15657 8076 15691
rect 8024 15648 8076 15657
rect 8300 15648 8352 15700
rect 11612 15691 11664 15700
rect 11612 15657 11621 15691
rect 11621 15657 11655 15691
rect 11655 15657 11664 15691
rect 11612 15648 11664 15657
rect 13728 15648 13780 15700
rect 21824 15648 21876 15700
rect 6460 15580 6512 15632
rect 7196 15580 7248 15632
rect 3148 15512 3200 15564
rect 2964 15487 3016 15496
rect 2964 15453 2973 15487
rect 2973 15453 3007 15487
rect 3007 15453 3016 15487
rect 2964 15444 3016 15453
rect 3884 15555 3936 15564
rect 3884 15521 3893 15555
rect 3893 15521 3927 15555
rect 3927 15521 3936 15555
rect 3884 15512 3936 15521
rect 3976 15555 4028 15564
rect 3976 15521 3985 15555
rect 3985 15521 4019 15555
rect 4019 15521 4028 15555
rect 3976 15512 4028 15521
rect 4712 15512 4764 15564
rect 7748 15555 7800 15564
rect 7748 15521 7757 15555
rect 7757 15521 7791 15555
rect 7791 15521 7800 15555
rect 7748 15512 7800 15521
rect 8208 15512 8260 15564
rect 8116 15444 8168 15496
rect 11336 15555 11388 15564
rect 11336 15521 11345 15555
rect 11345 15521 11379 15555
rect 11379 15521 11388 15555
rect 11336 15512 11388 15521
rect 10968 15487 11020 15496
rect 10968 15453 10977 15487
rect 10977 15453 11011 15487
rect 11011 15453 11020 15487
rect 10968 15444 11020 15453
rect 11244 15487 11296 15496
rect 11244 15453 11253 15487
rect 11253 15453 11287 15487
rect 11287 15453 11296 15487
rect 13268 15555 13320 15564
rect 13268 15521 13277 15555
rect 13277 15521 13311 15555
rect 13311 15521 13320 15555
rect 13268 15512 13320 15521
rect 13452 15512 13504 15564
rect 13820 15512 13872 15564
rect 11244 15444 11296 15453
rect 13360 15487 13412 15496
rect 13360 15453 13369 15487
rect 13369 15453 13403 15487
rect 13403 15453 13412 15487
rect 13360 15444 13412 15453
rect 4712 15376 4764 15428
rect 6368 15376 6420 15428
rect 8668 15376 8720 15428
rect 12900 15419 12952 15428
rect 12900 15385 12909 15419
rect 12909 15385 12943 15419
rect 12943 15385 12952 15419
rect 12900 15376 12952 15385
rect 15016 15555 15068 15564
rect 15016 15521 15025 15555
rect 15025 15521 15059 15555
rect 15059 15521 15068 15555
rect 15016 15512 15068 15521
rect 15200 15555 15252 15564
rect 15200 15521 15209 15555
rect 15209 15521 15243 15555
rect 15243 15521 15252 15555
rect 15200 15512 15252 15521
rect 15384 15512 15436 15564
rect 14924 15444 14976 15496
rect 21548 15580 21600 15632
rect 18512 15555 18564 15564
rect 18512 15521 18546 15555
rect 18546 15521 18564 15555
rect 18512 15512 18564 15521
rect 21088 15512 21140 15564
rect 22008 15512 22060 15564
rect 4252 15308 4304 15360
rect 8760 15308 8812 15360
rect 18236 15487 18288 15496
rect 18236 15453 18245 15487
rect 18245 15453 18279 15487
rect 18279 15453 18288 15487
rect 18236 15444 18288 15453
rect 21824 15487 21876 15496
rect 21824 15453 21833 15487
rect 21833 15453 21867 15487
rect 21867 15453 21876 15487
rect 21824 15444 21876 15453
rect 15936 15376 15988 15428
rect 21456 15376 21508 15428
rect 22468 15376 22520 15428
rect 15660 15351 15712 15360
rect 15660 15317 15669 15351
rect 15669 15317 15703 15351
rect 15703 15317 15712 15351
rect 15660 15308 15712 15317
rect 15752 15351 15804 15360
rect 15752 15317 15761 15351
rect 15761 15317 15795 15351
rect 15795 15317 15804 15351
rect 15752 15308 15804 15317
rect 19432 15308 19484 15360
rect 22284 15351 22336 15360
rect 22284 15317 22293 15351
rect 22293 15317 22327 15351
rect 22327 15317 22336 15351
rect 22284 15308 22336 15317
rect 3662 15206 3714 15258
rect 3726 15206 3778 15258
rect 3790 15206 3842 15258
rect 3854 15206 3906 15258
rect 3918 15206 3970 15258
rect 11244 15104 11296 15156
rect 13820 15104 13872 15156
rect 16028 15104 16080 15156
rect 17960 15104 18012 15156
rect 4252 15011 4304 15020
rect 4252 14977 4261 15011
rect 4261 14977 4295 15011
rect 4295 14977 4304 15011
rect 4252 14968 4304 14977
rect 4712 15011 4764 15020
rect 4712 14977 4721 15011
rect 4721 14977 4755 15011
rect 4755 14977 4764 15011
rect 4712 14968 4764 14977
rect 10968 15036 11020 15088
rect 16488 15036 16540 15088
rect 5908 14968 5960 15020
rect 15752 14968 15804 15020
rect 4160 14943 4212 14952
rect 4160 14909 4169 14943
rect 4169 14909 4203 14943
rect 4203 14909 4212 14943
rect 4160 14900 4212 14909
rect 4988 14900 5040 14952
rect 7012 14900 7064 14952
rect 11060 14900 11112 14952
rect 12624 14943 12676 14952
rect 12624 14909 12633 14943
rect 12633 14909 12667 14943
rect 12667 14909 12676 14943
rect 12624 14900 12676 14909
rect 14188 14900 14240 14952
rect 15476 14900 15528 14952
rect 16028 14943 16080 14952
rect 16028 14909 16037 14943
rect 16037 14909 16071 14943
rect 16071 14909 16080 14943
rect 16028 14900 16080 14909
rect 16580 14943 16632 14952
rect 16580 14909 16589 14943
rect 16589 14909 16623 14943
rect 16623 14909 16632 14943
rect 16580 14900 16632 14909
rect 16764 14943 16816 14952
rect 16764 14909 16773 14943
rect 16773 14909 16807 14943
rect 16807 14909 16816 14943
rect 16764 14900 16816 14909
rect 18420 15104 18472 15156
rect 21548 15104 21600 15156
rect 20352 14968 20404 15020
rect 20904 14968 20956 15020
rect 21456 14968 21508 15020
rect 19432 14900 19484 14952
rect 21364 14900 21416 14952
rect 22008 14943 22060 14952
rect 22008 14909 22017 14943
rect 22017 14909 22051 14943
rect 22051 14909 22060 14943
rect 22008 14900 22060 14909
rect 19892 14875 19944 14884
rect 19892 14841 19901 14875
rect 19901 14841 19935 14875
rect 19935 14841 19944 14875
rect 19892 14832 19944 14841
rect 20076 14875 20128 14884
rect 20076 14841 20085 14875
rect 20085 14841 20119 14875
rect 20119 14841 20128 14875
rect 20076 14832 20128 14841
rect 20628 14832 20680 14884
rect 21824 14875 21876 14884
rect 21824 14841 21833 14875
rect 21833 14841 21867 14875
rect 21867 14841 21876 14875
rect 21824 14832 21876 14841
rect 22560 14832 22612 14884
rect 22836 14832 22888 14884
rect 5172 14807 5224 14816
rect 5172 14773 5181 14807
rect 5181 14773 5215 14807
rect 5215 14773 5224 14807
rect 5172 14764 5224 14773
rect 5356 14807 5408 14816
rect 5356 14773 5365 14807
rect 5365 14773 5399 14807
rect 5399 14773 5408 14807
rect 5356 14764 5408 14773
rect 11520 14764 11572 14816
rect 12808 14764 12860 14816
rect 16396 14764 16448 14816
rect 4322 14662 4374 14714
rect 4386 14662 4438 14714
rect 4450 14662 4502 14714
rect 4514 14662 4566 14714
rect 4578 14662 4630 14714
rect 2964 14560 3016 14612
rect 3424 14560 3476 14612
rect 5356 14560 5408 14612
rect 4160 14492 4212 14544
rect 2780 14424 2832 14476
rect 2872 14467 2924 14476
rect 2872 14433 2881 14467
rect 2881 14433 2915 14467
rect 2915 14433 2924 14467
rect 2872 14424 2924 14433
rect 4252 14424 4304 14476
rect 5172 14467 5224 14476
rect 5172 14433 5181 14467
rect 5181 14433 5215 14467
rect 5215 14433 5224 14467
rect 5172 14424 5224 14433
rect 6092 14424 6144 14476
rect 7196 14424 7248 14476
rect 8024 14467 8076 14476
rect 8024 14433 8033 14467
rect 8033 14433 8067 14467
rect 8067 14433 8076 14467
rect 8024 14424 8076 14433
rect 9036 14424 9088 14476
rect 10048 14492 10100 14544
rect 15752 14535 15804 14544
rect 15752 14501 15761 14535
rect 15761 14501 15795 14535
rect 15795 14501 15804 14535
rect 15752 14492 15804 14501
rect 5448 14356 5500 14408
rect 5908 14399 5960 14408
rect 5908 14365 5917 14399
rect 5917 14365 5951 14399
rect 5951 14365 5960 14399
rect 5908 14356 5960 14365
rect 8392 14356 8444 14408
rect 15476 14424 15528 14476
rect 15660 14467 15712 14476
rect 15660 14433 15669 14467
rect 15669 14433 15703 14467
rect 15703 14433 15712 14467
rect 15660 14424 15712 14433
rect 15936 14467 15988 14476
rect 15936 14433 15945 14467
rect 15945 14433 15979 14467
rect 15979 14433 15988 14467
rect 15936 14424 15988 14433
rect 16396 14467 16448 14476
rect 16396 14433 16405 14467
rect 16405 14433 16439 14467
rect 16439 14433 16448 14467
rect 16396 14424 16448 14433
rect 16488 14467 16540 14476
rect 16488 14433 16497 14467
rect 16497 14433 16531 14467
rect 16531 14433 16540 14467
rect 16488 14424 16540 14433
rect 6000 14288 6052 14340
rect 17500 14356 17552 14408
rect 9680 14288 9732 14340
rect 15016 14288 15068 14340
rect 19340 14560 19392 14612
rect 17776 14424 17828 14476
rect 19432 14467 19484 14476
rect 19432 14433 19441 14467
rect 19441 14433 19475 14467
rect 19475 14433 19484 14467
rect 19432 14424 19484 14433
rect 19892 14424 19944 14476
rect 21088 14560 21140 14612
rect 19248 14356 19300 14408
rect 20352 14467 20404 14476
rect 20352 14433 20361 14467
rect 20361 14433 20395 14467
rect 20395 14433 20404 14467
rect 20352 14424 20404 14433
rect 20628 14424 20680 14476
rect 6736 14220 6788 14272
rect 8944 14220 8996 14272
rect 15384 14263 15436 14272
rect 15384 14229 15393 14263
rect 15393 14229 15427 14263
rect 15427 14229 15436 14263
rect 15384 14220 15436 14229
rect 16856 14220 16908 14272
rect 19616 14220 19668 14272
rect 20168 14263 20220 14272
rect 20168 14229 20177 14263
rect 20177 14229 20211 14263
rect 20211 14229 20220 14263
rect 20168 14220 20220 14229
rect 20812 14220 20864 14272
rect 3662 14118 3714 14170
rect 3726 14118 3778 14170
rect 3790 14118 3842 14170
rect 3854 14118 3906 14170
rect 3918 14118 3970 14170
rect 2780 13855 2832 13864
rect 2780 13821 2789 13855
rect 2789 13821 2823 13855
rect 2823 13821 2832 13855
rect 2780 13812 2832 13821
rect 2872 13855 2924 13864
rect 2872 13821 2881 13855
rect 2881 13821 2915 13855
rect 2915 13821 2924 13855
rect 2872 13812 2924 13821
rect 5172 13948 5224 14000
rect 3148 13880 3200 13932
rect 3424 13855 3476 13864
rect 3424 13821 3433 13855
rect 3433 13821 3467 13855
rect 3467 13821 3476 13855
rect 3424 13812 3476 13821
rect 5448 13880 5500 13932
rect 6000 13923 6052 13932
rect 6000 13889 6009 13923
rect 6009 13889 6043 13923
rect 6043 13889 6052 13923
rect 6000 13880 6052 13889
rect 6644 13923 6696 13932
rect 6644 13889 6653 13923
rect 6653 13889 6687 13923
rect 6687 13889 6696 13923
rect 6644 13880 6696 13889
rect 6092 13855 6144 13864
rect 6092 13821 6101 13855
rect 6101 13821 6135 13855
rect 6135 13821 6144 13855
rect 6092 13812 6144 13821
rect 6736 13855 6788 13864
rect 6736 13821 6745 13855
rect 6745 13821 6779 13855
rect 6779 13821 6788 13855
rect 6736 13812 6788 13821
rect 3148 13744 3200 13796
rect 3516 13787 3568 13796
rect 3516 13753 3525 13787
rect 3525 13753 3559 13787
rect 3559 13753 3568 13787
rect 3516 13744 3568 13753
rect 6644 13744 6696 13796
rect 9496 14016 9548 14068
rect 11244 14016 11296 14068
rect 13912 14016 13964 14068
rect 15660 14016 15712 14068
rect 16212 14016 16264 14068
rect 17500 14016 17552 14068
rect 20168 14059 20220 14068
rect 20168 14025 20177 14059
rect 20177 14025 20211 14059
rect 20211 14025 20220 14059
rect 20168 14016 20220 14025
rect 8852 13948 8904 14000
rect 8024 13855 8076 13864
rect 8024 13821 8063 13855
rect 8063 13821 8076 13855
rect 8024 13812 8076 13821
rect 8392 13812 8444 13864
rect 8944 13923 8996 13932
rect 8944 13889 8953 13923
rect 8953 13889 8987 13923
rect 8987 13889 8996 13923
rect 8944 13880 8996 13889
rect 8852 13744 8904 13796
rect 9036 13855 9088 13864
rect 9036 13821 9045 13855
rect 9045 13821 9079 13855
rect 9079 13821 9088 13855
rect 9036 13812 9088 13821
rect 11060 13812 11112 13864
rect 11244 13855 11296 13864
rect 11244 13821 11253 13855
rect 11253 13821 11287 13855
rect 11287 13821 11296 13855
rect 11244 13812 11296 13821
rect 17776 13948 17828 14000
rect 13268 13880 13320 13932
rect 11520 13855 11572 13864
rect 11520 13821 11529 13855
rect 11529 13821 11563 13855
rect 11563 13821 11572 13855
rect 11520 13812 11572 13821
rect 12900 13812 12952 13864
rect 13636 13855 13688 13864
rect 13636 13821 13645 13855
rect 13645 13821 13679 13855
rect 13679 13821 13688 13855
rect 13636 13812 13688 13821
rect 3792 13719 3844 13728
rect 3792 13685 3801 13719
rect 3801 13685 3835 13719
rect 3835 13685 3844 13719
rect 3792 13676 3844 13685
rect 5724 13719 5776 13728
rect 5724 13685 5733 13719
rect 5733 13685 5767 13719
rect 5767 13685 5776 13719
rect 5724 13676 5776 13685
rect 8668 13719 8720 13728
rect 8668 13685 8677 13719
rect 8677 13685 8711 13719
rect 8711 13685 8720 13719
rect 8668 13676 8720 13685
rect 10232 13676 10284 13728
rect 12348 13744 12400 13796
rect 14556 13812 14608 13864
rect 15384 13812 15436 13864
rect 16856 13812 16908 13864
rect 18236 13880 18288 13932
rect 18512 13880 18564 13932
rect 20904 14059 20956 14068
rect 20904 14025 20913 14059
rect 20913 14025 20947 14059
rect 20947 14025 20956 14059
rect 20904 14016 20956 14025
rect 22008 14016 22060 14068
rect 19432 13880 19484 13932
rect 19616 13923 19668 13932
rect 19616 13889 19625 13923
rect 19625 13889 19659 13923
rect 19659 13889 19668 13923
rect 19616 13880 19668 13889
rect 19340 13812 19392 13864
rect 21456 13923 21508 13932
rect 21456 13889 21465 13923
rect 21465 13889 21499 13923
rect 21499 13889 21508 13923
rect 21456 13880 21508 13889
rect 20812 13812 20864 13864
rect 20168 13787 20220 13796
rect 20168 13753 20177 13787
rect 20177 13753 20211 13787
rect 20211 13753 20220 13787
rect 20168 13744 20220 13753
rect 21548 13855 21600 13864
rect 21548 13821 21557 13855
rect 21557 13821 21591 13855
rect 21591 13821 21600 13855
rect 21548 13812 21600 13821
rect 21088 13787 21140 13796
rect 21088 13753 21097 13787
rect 21097 13753 21131 13787
rect 21131 13753 21140 13787
rect 21088 13744 21140 13753
rect 22468 13855 22520 13864
rect 22468 13821 22477 13855
rect 22477 13821 22511 13855
rect 22511 13821 22520 13855
rect 22468 13812 22520 13821
rect 22560 13744 22612 13796
rect 12716 13676 12768 13728
rect 20720 13676 20772 13728
rect 4322 13574 4374 13626
rect 4386 13574 4438 13626
rect 4450 13574 4502 13626
rect 4514 13574 4566 13626
rect 4578 13574 4630 13626
rect 3792 13404 3844 13456
rect 5724 13404 5776 13456
rect 9496 13447 9548 13456
rect 9496 13413 9505 13447
rect 9505 13413 9539 13447
rect 9539 13413 9548 13447
rect 9496 13404 9548 13413
rect 12900 13472 12952 13524
rect 6000 13379 6052 13388
rect 6000 13345 6009 13379
rect 6009 13345 6043 13379
rect 6043 13345 6052 13379
rect 6000 13336 6052 13345
rect 7012 13336 7064 13388
rect 8208 13336 8260 13388
rect 4712 13268 4764 13320
rect 9680 13268 9732 13320
rect 10232 13379 10284 13388
rect 10232 13345 10241 13379
rect 10241 13345 10275 13379
rect 10275 13345 10284 13379
rect 10232 13336 10284 13345
rect 6644 13200 6696 13252
rect 9956 13200 10008 13252
rect 12348 13336 12400 13388
rect 12716 13379 12768 13388
rect 12716 13345 12725 13379
rect 12725 13345 12759 13379
rect 12759 13345 12768 13379
rect 12716 13336 12768 13345
rect 12808 13379 12860 13388
rect 12808 13345 12817 13379
rect 12817 13345 12851 13379
rect 12851 13345 12860 13379
rect 12808 13336 12860 13345
rect 12900 13379 12952 13388
rect 12900 13345 12909 13379
rect 12909 13345 12943 13379
rect 12943 13345 12952 13379
rect 12900 13336 12952 13345
rect 13176 13379 13228 13388
rect 13176 13345 13185 13379
rect 13185 13345 13219 13379
rect 13219 13345 13228 13379
rect 13176 13336 13228 13345
rect 13268 13379 13320 13388
rect 13268 13345 13277 13379
rect 13277 13345 13311 13379
rect 13311 13345 13320 13379
rect 13268 13336 13320 13345
rect 13636 13404 13688 13456
rect 13820 13472 13872 13524
rect 17500 13447 17552 13456
rect 17500 13413 17509 13447
rect 17509 13413 17543 13447
rect 17543 13413 17552 13447
rect 17500 13404 17552 13413
rect 12348 13200 12400 13252
rect 17224 13336 17276 13388
rect 21456 13379 21508 13388
rect 21456 13345 21465 13379
rect 21465 13345 21499 13379
rect 21499 13345 21508 13379
rect 21456 13336 21508 13345
rect 3424 13132 3476 13184
rect 9680 13175 9732 13184
rect 9680 13141 9689 13175
rect 9689 13141 9723 13175
rect 9723 13141 9732 13175
rect 9680 13132 9732 13141
rect 10416 13175 10468 13184
rect 10416 13141 10425 13175
rect 10425 13141 10459 13175
rect 10459 13141 10468 13175
rect 10416 13132 10468 13141
rect 10508 13175 10560 13184
rect 10508 13141 10517 13175
rect 10517 13141 10551 13175
rect 10551 13141 10560 13175
rect 10508 13132 10560 13141
rect 13360 13132 13412 13184
rect 13820 13175 13872 13184
rect 13820 13141 13829 13175
rect 13829 13141 13863 13175
rect 13863 13141 13872 13175
rect 13820 13132 13872 13141
rect 17316 13200 17368 13252
rect 19064 13200 19116 13252
rect 21916 13472 21968 13524
rect 21732 13404 21784 13456
rect 22284 13404 22336 13456
rect 21732 13311 21784 13320
rect 21732 13277 21741 13311
rect 21741 13277 21775 13311
rect 21775 13277 21784 13311
rect 21732 13268 21784 13277
rect 22468 13379 22520 13388
rect 22468 13345 22477 13379
rect 22477 13345 22511 13379
rect 22511 13345 22520 13379
rect 22468 13336 22520 13345
rect 22192 13200 22244 13252
rect 22836 13311 22888 13320
rect 22836 13277 22845 13311
rect 22845 13277 22879 13311
rect 22879 13277 22888 13311
rect 22836 13268 22888 13277
rect 14280 13175 14332 13184
rect 14280 13141 14289 13175
rect 14289 13141 14323 13175
rect 14323 13141 14332 13175
rect 14280 13132 14332 13141
rect 17776 13132 17828 13184
rect 22008 13132 22060 13184
rect 3662 13030 3714 13082
rect 3726 13030 3778 13082
rect 3790 13030 3842 13082
rect 3854 13030 3906 13082
rect 3918 13030 3970 13082
rect 8760 12971 8812 12980
rect 8760 12937 8769 12971
rect 8769 12937 8803 12971
rect 8803 12937 8812 12971
rect 8760 12928 8812 12937
rect 9404 12928 9456 12980
rect 5264 12792 5316 12844
rect 6920 12835 6972 12844
rect 6920 12801 6929 12835
rect 6929 12801 6963 12835
rect 6963 12801 6972 12835
rect 6920 12792 6972 12801
rect 7196 12835 7248 12844
rect 7196 12801 7205 12835
rect 7205 12801 7239 12835
rect 7239 12801 7248 12835
rect 7196 12792 7248 12801
rect 4988 12724 5040 12776
rect 5356 12724 5408 12776
rect 9680 12860 9732 12912
rect 8576 12792 8628 12844
rect 8668 12724 8720 12776
rect 8852 12724 8904 12776
rect 10416 12792 10468 12844
rect 12440 12928 12492 12980
rect 12532 12928 12584 12980
rect 13268 12928 13320 12980
rect 14280 12928 14332 12980
rect 17776 12928 17828 12980
rect 18328 12928 18380 12980
rect 20168 12928 20220 12980
rect 21732 12971 21784 12980
rect 21732 12937 21741 12971
rect 21741 12937 21775 12971
rect 21775 12937 21784 12971
rect 21732 12928 21784 12937
rect 12256 12792 12308 12844
rect 19524 12860 19576 12912
rect 21640 12860 21692 12912
rect 12808 12792 12860 12844
rect 8392 12656 8444 12708
rect 4252 12588 4304 12640
rect 4804 12588 4856 12640
rect 7932 12588 7984 12640
rect 9404 12767 9456 12776
rect 9404 12733 9413 12767
rect 9413 12733 9447 12767
rect 9447 12733 9456 12767
rect 9404 12724 9456 12733
rect 11888 12767 11940 12776
rect 11888 12733 11897 12767
rect 11897 12733 11931 12767
rect 11931 12733 11940 12767
rect 11888 12724 11940 12733
rect 10692 12656 10744 12708
rect 12440 12767 12492 12776
rect 12440 12733 12449 12767
rect 12449 12733 12483 12767
rect 12483 12733 12492 12767
rect 12440 12724 12492 12733
rect 12716 12724 12768 12776
rect 13452 12792 13504 12844
rect 13820 12767 13872 12776
rect 13820 12733 13829 12767
rect 13829 12733 13863 12767
rect 13863 12733 13872 12767
rect 13820 12724 13872 12733
rect 15292 12792 15344 12844
rect 17316 12792 17368 12844
rect 17224 12767 17276 12776
rect 17224 12733 17233 12767
rect 17233 12733 17267 12767
rect 17267 12733 17276 12767
rect 17224 12724 17276 12733
rect 17500 12792 17552 12844
rect 18052 12835 18104 12844
rect 18052 12801 18061 12835
rect 18061 12801 18095 12835
rect 18095 12801 18104 12835
rect 18052 12792 18104 12801
rect 21824 12792 21876 12844
rect 9404 12631 9456 12640
rect 9404 12597 9413 12631
rect 9413 12597 9447 12631
rect 9447 12597 9456 12631
rect 9404 12588 9456 12597
rect 11704 12631 11756 12640
rect 11704 12597 11713 12631
rect 11713 12597 11747 12631
rect 11747 12597 11756 12631
rect 11704 12588 11756 12597
rect 11888 12588 11940 12640
rect 12440 12588 12492 12640
rect 15936 12656 15988 12708
rect 18144 12724 18196 12776
rect 18236 12767 18288 12776
rect 18236 12733 18245 12767
rect 18245 12733 18279 12767
rect 18279 12733 18288 12767
rect 18236 12724 18288 12733
rect 17960 12699 18012 12708
rect 17960 12665 17969 12699
rect 17969 12665 18003 12699
rect 18003 12665 18012 12699
rect 17960 12656 18012 12665
rect 13268 12631 13320 12640
rect 13268 12597 13277 12631
rect 13277 12597 13311 12631
rect 13311 12597 13320 12631
rect 13268 12588 13320 12597
rect 14372 12588 14424 12640
rect 14924 12631 14976 12640
rect 14924 12597 14933 12631
rect 14933 12597 14967 12631
rect 14967 12597 14976 12631
rect 14924 12588 14976 12597
rect 17684 12631 17736 12640
rect 17684 12597 17709 12631
rect 17709 12597 17736 12631
rect 17684 12588 17736 12597
rect 18880 12588 18932 12640
rect 22468 12656 22520 12708
rect 22192 12588 22244 12640
rect 4322 12486 4374 12538
rect 4386 12486 4438 12538
rect 4450 12486 4502 12538
rect 4514 12486 4566 12538
rect 4578 12486 4630 12538
rect 2780 12384 2832 12436
rect 5356 12427 5408 12436
rect 5356 12393 5365 12427
rect 5365 12393 5399 12427
rect 5399 12393 5408 12427
rect 5356 12384 5408 12393
rect 9404 12384 9456 12436
rect 4252 12359 4304 12368
rect 4252 12325 4286 12359
rect 4286 12325 4304 12359
rect 4252 12316 4304 12325
rect 8576 12316 8628 12368
rect 8852 12359 8904 12368
rect 8852 12325 8861 12359
rect 8861 12325 8895 12359
rect 8895 12325 8904 12359
rect 8852 12316 8904 12325
rect 9680 12359 9732 12368
rect 9680 12325 9689 12359
rect 9689 12325 9723 12359
rect 9723 12325 9732 12359
rect 9680 12316 9732 12325
rect 4620 12248 4672 12300
rect 7196 12248 7248 12300
rect 7380 12248 7432 12300
rect 3240 12223 3292 12232
rect 3240 12189 3249 12223
rect 3249 12189 3283 12223
rect 3283 12189 3292 12223
rect 3240 12180 3292 12189
rect 3332 12223 3384 12232
rect 3332 12189 3341 12223
rect 3341 12189 3375 12223
rect 3375 12189 3384 12223
rect 3332 12180 3384 12189
rect 7840 12180 7892 12232
rect 8208 12291 8260 12300
rect 8208 12257 8217 12291
rect 8217 12257 8251 12291
rect 8251 12257 8260 12291
rect 8208 12248 8260 12257
rect 8760 12248 8812 12300
rect 9956 12291 10008 12300
rect 9956 12257 9965 12291
rect 9965 12257 9999 12291
rect 9999 12257 10008 12291
rect 9956 12248 10008 12257
rect 10232 12248 10284 12300
rect 10508 12248 10560 12300
rect 12440 12427 12492 12436
rect 12440 12393 12449 12427
rect 12449 12393 12483 12427
rect 12483 12393 12492 12427
rect 12440 12384 12492 12393
rect 14924 12316 14976 12368
rect 16672 12359 16724 12368
rect 16672 12325 16681 12359
rect 16681 12325 16715 12359
rect 16715 12325 16724 12359
rect 16672 12316 16724 12325
rect 17776 12427 17828 12436
rect 17776 12393 17785 12427
rect 17785 12393 17819 12427
rect 17819 12393 17828 12427
rect 17776 12384 17828 12393
rect 18236 12384 18288 12436
rect 18328 12384 18380 12436
rect 22744 12384 22796 12436
rect 18144 12316 18196 12368
rect 18880 12359 18932 12368
rect 18880 12325 18889 12359
rect 18889 12325 18923 12359
rect 18923 12325 18932 12359
rect 18880 12316 18932 12325
rect 12348 12291 12400 12300
rect 12348 12257 12357 12291
rect 12357 12257 12391 12291
rect 12391 12257 12400 12291
rect 12348 12248 12400 12257
rect 12532 12291 12584 12300
rect 12532 12257 12541 12291
rect 12541 12257 12575 12291
rect 12575 12257 12584 12291
rect 12532 12248 12584 12257
rect 13268 12291 13320 12300
rect 13268 12257 13277 12291
rect 13277 12257 13311 12291
rect 13311 12257 13320 12291
rect 13268 12248 13320 12257
rect 13360 12291 13412 12300
rect 13360 12257 13369 12291
rect 13369 12257 13403 12291
rect 13403 12257 13412 12291
rect 13360 12248 13412 12257
rect 13452 12291 13504 12300
rect 13452 12257 13461 12291
rect 13461 12257 13495 12291
rect 13495 12257 13504 12291
rect 13452 12248 13504 12257
rect 14280 12248 14332 12300
rect 17132 12291 17184 12300
rect 17132 12257 17141 12291
rect 17141 12257 17175 12291
rect 17175 12257 17184 12291
rect 17132 12248 17184 12257
rect 17224 12291 17276 12300
rect 17224 12257 17233 12291
rect 17233 12257 17267 12291
rect 17267 12257 17276 12291
rect 17224 12248 17276 12257
rect 17684 12291 17736 12300
rect 17684 12257 17693 12291
rect 17693 12257 17727 12291
rect 17727 12257 17736 12291
rect 17684 12248 17736 12257
rect 18420 12291 18472 12300
rect 18420 12257 18429 12291
rect 18429 12257 18463 12291
rect 18463 12257 18472 12291
rect 18420 12248 18472 12257
rect 13544 12223 13596 12232
rect 13544 12189 13553 12223
rect 13553 12189 13587 12223
rect 13587 12189 13596 12223
rect 13544 12180 13596 12189
rect 14556 12223 14608 12232
rect 14556 12189 14565 12223
rect 14565 12189 14599 12223
rect 14599 12189 14608 12223
rect 14556 12180 14608 12189
rect 10692 12112 10744 12164
rect 4344 12044 4396 12096
rect 8392 12044 8444 12096
rect 9312 12044 9364 12096
rect 9680 12044 9732 12096
rect 10508 12087 10560 12096
rect 10508 12053 10517 12087
rect 10517 12053 10551 12087
rect 10551 12053 10560 12087
rect 10508 12044 10560 12053
rect 13084 12087 13136 12096
rect 13084 12053 13093 12087
rect 13093 12053 13127 12087
rect 13127 12053 13136 12087
rect 13084 12044 13136 12053
rect 18512 12223 18564 12232
rect 18512 12189 18521 12223
rect 18521 12189 18555 12223
rect 18555 12189 18564 12223
rect 18512 12180 18564 12189
rect 14924 12044 14976 12096
rect 15936 12087 15988 12096
rect 15936 12053 15945 12087
rect 15945 12053 15979 12087
rect 15979 12053 15988 12087
rect 15936 12044 15988 12053
rect 16120 12044 16172 12096
rect 16580 12044 16632 12096
rect 20352 12316 20404 12368
rect 21548 12248 21600 12300
rect 21916 12248 21968 12300
rect 22100 12248 22152 12300
rect 23020 12291 23072 12300
rect 23020 12257 23029 12291
rect 23029 12257 23063 12291
rect 23063 12257 23072 12291
rect 23020 12248 23072 12257
rect 20996 12180 21048 12232
rect 21548 12112 21600 12164
rect 17040 12087 17092 12096
rect 17040 12053 17049 12087
rect 17049 12053 17083 12087
rect 17083 12053 17092 12087
rect 17040 12044 17092 12053
rect 17316 12044 17368 12096
rect 19524 12044 19576 12096
rect 20720 12044 20772 12096
rect 22008 12087 22060 12096
rect 22008 12053 22017 12087
rect 22017 12053 22051 12087
rect 22051 12053 22060 12087
rect 22008 12044 22060 12053
rect 3662 11942 3714 11994
rect 3726 11942 3778 11994
rect 3790 11942 3842 11994
rect 3854 11942 3906 11994
rect 3918 11942 3970 11994
rect 3332 11840 3384 11892
rect 10232 11840 10284 11892
rect 16212 11883 16264 11892
rect 16212 11849 16221 11883
rect 16221 11849 16255 11883
rect 16255 11849 16264 11883
rect 16212 11840 16264 11849
rect 16580 11840 16632 11892
rect 17132 11840 17184 11892
rect 18052 11840 18104 11892
rect 19524 11883 19576 11892
rect 19524 11849 19533 11883
rect 19533 11849 19567 11883
rect 19567 11849 19576 11883
rect 19524 11840 19576 11849
rect 20352 11840 20404 11892
rect 4620 11747 4672 11756
rect 4620 11713 4629 11747
rect 4629 11713 4663 11747
rect 4663 11713 4672 11747
rect 4620 11704 4672 11713
rect 4896 11704 4948 11756
rect 5264 11747 5316 11756
rect 5264 11713 5273 11747
rect 5273 11713 5307 11747
rect 5307 11713 5316 11747
rect 5264 11704 5316 11713
rect 7564 11772 7616 11824
rect 9864 11704 9916 11756
rect 10508 11704 10560 11756
rect 10692 11747 10744 11756
rect 10692 11713 10701 11747
rect 10701 11713 10735 11747
rect 10735 11713 10744 11747
rect 10692 11704 10744 11713
rect 14924 11747 14976 11756
rect 14924 11713 14933 11747
rect 14933 11713 14967 11747
rect 14967 11713 14976 11747
rect 14924 11704 14976 11713
rect 20812 11840 20864 11892
rect 21180 11840 21232 11892
rect 17040 11704 17092 11756
rect 4344 11679 4396 11688
rect 4344 11645 4362 11679
rect 4362 11645 4396 11679
rect 4344 11636 4396 11645
rect 7196 11679 7248 11688
rect 7196 11645 7205 11679
rect 7205 11645 7239 11679
rect 7239 11645 7248 11679
rect 7196 11636 7248 11645
rect 7380 11636 7432 11688
rect 7932 11679 7984 11688
rect 7932 11645 7941 11679
rect 7941 11645 7975 11679
rect 7975 11645 7984 11679
rect 7932 11636 7984 11645
rect 8392 11679 8444 11688
rect 8392 11645 8401 11679
rect 8401 11645 8435 11679
rect 8435 11645 8444 11679
rect 8392 11636 8444 11645
rect 9312 11679 9364 11688
rect 9312 11645 9321 11679
rect 9321 11645 9355 11679
rect 9355 11645 9364 11679
rect 9312 11636 9364 11645
rect 9404 11679 9456 11688
rect 9404 11645 9413 11679
rect 9413 11645 9447 11679
rect 9447 11645 9456 11679
rect 9404 11636 9456 11645
rect 9956 11636 10008 11688
rect 3240 11568 3292 11620
rect 7012 11611 7064 11620
rect 7012 11577 7021 11611
rect 7021 11577 7055 11611
rect 7055 11577 7064 11611
rect 7012 11568 7064 11577
rect 10692 11568 10744 11620
rect 10876 11679 10928 11688
rect 10876 11645 10885 11679
rect 10885 11645 10919 11679
rect 10919 11645 10928 11679
rect 10876 11636 10928 11645
rect 13084 11636 13136 11688
rect 15660 11636 15712 11688
rect 15016 11568 15068 11620
rect 16120 11679 16172 11688
rect 16120 11645 16129 11679
rect 16129 11645 16163 11679
rect 16163 11645 16172 11679
rect 16120 11636 16172 11645
rect 17316 11679 17368 11688
rect 17316 11645 17325 11679
rect 17325 11645 17359 11679
rect 17359 11645 17368 11679
rect 17316 11636 17368 11645
rect 21640 11883 21692 11892
rect 21640 11849 21649 11883
rect 21649 11849 21683 11883
rect 21683 11849 21692 11883
rect 21640 11840 21692 11849
rect 20720 11636 20772 11688
rect 22376 11636 22428 11688
rect 19524 11568 19576 11620
rect 21824 11568 21876 11620
rect 4712 11543 4764 11552
rect 4712 11509 4721 11543
rect 4721 11509 4755 11543
rect 4755 11509 4764 11543
rect 4712 11500 4764 11509
rect 5080 11543 5132 11552
rect 5080 11509 5089 11543
rect 5089 11509 5123 11543
rect 5123 11509 5132 11543
rect 5080 11500 5132 11509
rect 8024 11543 8076 11552
rect 8024 11509 8033 11543
rect 8033 11509 8067 11543
rect 8067 11509 8076 11543
rect 8024 11500 8076 11509
rect 8760 11543 8812 11552
rect 8760 11509 8769 11543
rect 8769 11509 8803 11543
rect 8803 11509 8812 11543
rect 8760 11500 8812 11509
rect 9128 11543 9180 11552
rect 9128 11509 9137 11543
rect 9137 11509 9171 11543
rect 9171 11509 9180 11543
rect 9128 11500 9180 11509
rect 10416 11543 10468 11552
rect 10416 11509 10425 11543
rect 10425 11509 10459 11543
rect 10459 11509 10468 11543
rect 10416 11500 10468 11509
rect 13636 11500 13688 11552
rect 4322 11398 4374 11450
rect 4386 11398 4438 11450
rect 4450 11398 4502 11450
rect 4514 11398 4566 11450
rect 4578 11398 4630 11450
rect 5080 11296 5132 11348
rect 6184 11296 6236 11348
rect 10876 11296 10928 11348
rect 4712 11228 4764 11280
rect 7012 11228 7064 11280
rect 12256 11296 12308 11348
rect 13544 11339 13596 11348
rect 13544 11305 13553 11339
rect 13553 11305 13587 11339
rect 13587 11305 13596 11339
rect 13544 11296 13596 11305
rect 18052 11296 18104 11348
rect 21824 11339 21876 11348
rect 21824 11305 21833 11339
rect 21833 11305 21867 11339
rect 21867 11305 21876 11339
rect 21824 11296 21876 11305
rect 6736 11160 6788 11212
rect 8024 11203 8076 11212
rect 8024 11169 8033 11203
rect 8033 11169 8067 11203
rect 8067 11169 8076 11203
rect 8024 11160 8076 11169
rect 8760 11160 8812 11212
rect 10508 11203 10560 11212
rect 10508 11169 10517 11203
rect 10517 11169 10551 11203
rect 10551 11169 10560 11203
rect 10508 11160 10560 11169
rect 18144 11228 18196 11280
rect 19340 11228 19392 11280
rect 20628 11228 20680 11280
rect 21548 11228 21600 11280
rect 22008 11271 22060 11280
rect 22008 11237 22017 11271
rect 22017 11237 22051 11271
rect 22051 11237 22060 11271
rect 22008 11228 22060 11237
rect 11244 11203 11296 11212
rect 11244 11169 11253 11203
rect 11253 11169 11287 11203
rect 11287 11169 11296 11203
rect 11244 11160 11296 11169
rect 11704 11203 11756 11212
rect 11704 11169 11713 11203
rect 11713 11169 11747 11203
rect 11747 11169 11756 11203
rect 11704 11160 11756 11169
rect 12440 11160 12492 11212
rect 15476 11160 15528 11212
rect 16120 11160 16172 11212
rect 19156 11160 19208 11212
rect 3240 11135 3292 11144
rect 3240 11101 3249 11135
rect 3249 11101 3283 11135
rect 3283 11101 3292 11135
rect 3240 11092 3292 11101
rect 5264 11092 5316 11144
rect 10692 11092 10744 11144
rect 12900 11092 12952 11144
rect 13636 11092 13688 11144
rect 15660 11135 15712 11144
rect 15660 11101 15669 11135
rect 15669 11101 15703 11135
rect 15703 11101 15712 11135
rect 15660 11092 15712 11101
rect 19340 11092 19392 11144
rect 20628 11135 20680 11144
rect 20628 11101 20637 11135
rect 20637 11101 20671 11135
rect 20671 11101 20680 11135
rect 20628 11092 20680 11101
rect 20720 11135 20772 11144
rect 20720 11101 20729 11135
rect 20729 11101 20763 11135
rect 20763 11101 20772 11135
rect 20720 11092 20772 11101
rect 20812 11024 20864 11076
rect 20904 11024 20956 11076
rect 22100 11024 22152 11076
rect 5632 10956 5684 11008
rect 8116 10999 8168 11008
rect 8116 10965 8125 10999
rect 8125 10965 8159 10999
rect 8159 10965 8168 10999
rect 8116 10956 8168 10965
rect 11612 10999 11664 11008
rect 11612 10965 11621 10999
rect 11621 10965 11655 10999
rect 11655 10965 11664 10999
rect 11612 10956 11664 10965
rect 15936 10999 15988 11008
rect 15936 10965 15945 10999
rect 15945 10965 15979 10999
rect 15979 10965 15988 10999
rect 15936 10956 15988 10965
rect 18420 10999 18472 11008
rect 18420 10965 18429 10999
rect 18429 10965 18463 10999
rect 18463 10965 18472 10999
rect 18420 10956 18472 10965
rect 19156 10956 19208 11008
rect 19524 10956 19576 11008
rect 19892 10956 19944 11008
rect 3662 10854 3714 10906
rect 3726 10854 3778 10906
rect 3790 10854 3842 10906
rect 3854 10854 3906 10906
rect 3918 10854 3970 10906
rect 6736 10795 6788 10804
rect 6736 10761 6745 10795
rect 6745 10761 6779 10795
rect 6779 10761 6788 10795
rect 6736 10752 6788 10761
rect 8116 10752 8168 10804
rect 10508 10752 10560 10804
rect 10968 10795 11020 10804
rect 10968 10761 10977 10795
rect 10977 10761 11011 10795
rect 11011 10761 11020 10795
rect 10968 10752 11020 10761
rect 11244 10752 11296 10804
rect 18512 10752 18564 10804
rect 19340 10795 19392 10804
rect 19340 10761 19349 10795
rect 19349 10761 19383 10795
rect 19383 10761 19392 10795
rect 19340 10752 19392 10761
rect 20812 10752 20864 10804
rect 21640 10752 21692 10804
rect 19156 10684 19208 10736
rect 20904 10684 20956 10736
rect 14096 10659 14148 10668
rect 14096 10625 14105 10659
rect 14105 10625 14139 10659
rect 14139 10625 14148 10659
rect 14096 10616 14148 10625
rect 14280 10659 14332 10668
rect 14280 10625 14289 10659
rect 14289 10625 14323 10659
rect 14323 10625 14332 10659
rect 14280 10616 14332 10625
rect 14556 10616 14608 10668
rect 5356 10591 5408 10600
rect 5356 10557 5365 10591
rect 5365 10557 5399 10591
rect 5399 10557 5408 10591
rect 5356 10548 5408 10557
rect 5632 10591 5684 10600
rect 5632 10557 5666 10591
rect 5666 10557 5684 10591
rect 5632 10548 5684 10557
rect 7012 10548 7064 10600
rect 7564 10591 7616 10600
rect 7564 10557 7573 10591
rect 7573 10557 7607 10591
rect 7607 10557 7616 10591
rect 7564 10548 7616 10557
rect 7840 10591 7892 10600
rect 7840 10557 7849 10591
rect 7849 10557 7883 10591
rect 7883 10557 7892 10591
rect 7840 10548 7892 10557
rect 7288 10523 7340 10532
rect 7288 10489 7297 10523
rect 7297 10489 7331 10523
rect 7331 10489 7340 10523
rect 7288 10480 7340 10489
rect 8116 10480 8168 10532
rect 8760 10548 8812 10600
rect 9128 10591 9180 10600
rect 9128 10557 9137 10591
rect 9137 10557 9171 10591
rect 9171 10557 9180 10591
rect 9128 10548 9180 10557
rect 9404 10480 9456 10532
rect 10416 10548 10468 10600
rect 11612 10548 11664 10600
rect 19248 10548 19300 10600
rect 21180 10548 21232 10600
rect 7012 10455 7064 10464
rect 7012 10421 7021 10455
rect 7021 10421 7055 10455
rect 7055 10421 7064 10455
rect 7012 10412 7064 10421
rect 8852 10412 8904 10464
rect 10508 10412 10560 10464
rect 13820 10412 13872 10464
rect 13912 10412 13964 10464
rect 18420 10412 18472 10464
rect 20076 10480 20128 10532
rect 20812 10523 20864 10532
rect 20812 10489 20821 10523
rect 20821 10489 20855 10523
rect 20855 10489 20864 10523
rect 20812 10480 20864 10489
rect 18880 10455 18932 10464
rect 18880 10421 18889 10455
rect 18889 10421 18923 10455
rect 18923 10421 18932 10455
rect 18880 10412 18932 10421
rect 19524 10412 19576 10464
rect 4322 10310 4374 10362
rect 4386 10310 4438 10362
rect 4450 10310 4502 10362
rect 4514 10310 4566 10362
rect 4578 10310 4630 10362
rect 5448 10208 5500 10260
rect 7288 10208 7340 10260
rect 7748 10208 7800 10260
rect 8116 10251 8168 10260
rect 8116 10217 8125 10251
rect 8125 10217 8159 10251
rect 8159 10217 8168 10251
rect 8116 10208 8168 10217
rect 3332 10115 3384 10124
rect 3332 10081 3341 10115
rect 3341 10081 3375 10115
rect 3375 10081 3384 10115
rect 3332 10072 3384 10081
rect 3516 10004 3568 10056
rect 7012 10140 7064 10192
rect 4896 10072 4948 10124
rect 5356 10072 5408 10124
rect 4712 10004 4764 10056
rect 5080 10047 5132 10056
rect 5080 10013 5089 10047
rect 5089 10013 5123 10047
rect 5123 10013 5132 10047
rect 5080 10004 5132 10013
rect 7840 10072 7892 10124
rect 14004 10072 14056 10124
rect 14372 10115 14424 10124
rect 14372 10081 14381 10115
rect 14381 10081 14415 10115
rect 14415 10081 14424 10115
rect 14372 10072 14424 10081
rect 14556 10115 14608 10124
rect 14556 10081 14565 10115
rect 14565 10081 14599 10115
rect 14599 10081 14608 10115
rect 14556 10072 14608 10081
rect 9404 10004 9456 10056
rect 15752 10183 15804 10192
rect 15752 10149 15777 10183
rect 15777 10149 15804 10183
rect 17960 10208 18012 10260
rect 18144 10251 18196 10260
rect 18144 10217 18153 10251
rect 18153 10217 18187 10251
rect 18187 10217 18196 10251
rect 18144 10208 18196 10217
rect 18512 10251 18564 10260
rect 18512 10217 18521 10251
rect 18521 10217 18555 10251
rect 18555 10217 18564 10251
rect 18512 10208 18564 10217
rect 20076 10251 20128 10260
rect 20076 10217 20085 10251
rect 20085 10217 20119 10251
rect 20119 10217 20128 10251
rect 20076 10208 20128 10217
rect 20904 10208 20956 10260
rect 15752 10140 15804 10149
rect 16580 10072 16632 10124
rect 16764 10115 16816 10124
rect 16764 10081 16773 10115
rect 16773 10081 16807 10115
rect 16807 10081 16816 10115
rect 16764 10072 16816 10081
rect 18880 10140 18932 10192
rect 20996 10140 21048 10192
rect 18052 10115 18104 10124
rect 18052 10081 18061 10115
rect 18061 10081 18095 10115
rect 18095 10081 18104 10115
rect 18052 10072 18104 10081
rect 18420 10072 18472 10124
rect 19524 10115 19576 10124
rect 19524 10081 19533 10115
rect 19533 10081 19567 10115
rect 19567 10081 19576 10115
rect 19524 10072 19576 10081
rect 20720 10072 20772 10124
rect 21548 10140 21600 10192
rect 22192 10140 22244 10192
rect 22468 10140 22520 10192
rect 22560 10183 22612 10192
rect 22560 10149 22569 10183
rect 22569 10149 22603 10183
rect 22603 10149 22612 10183
rect 22560 10140 22612 10149
rect 4068 9868 4120 9920
rect 4804 9936 4856 9988
rect 4620 9868 4672 9920
rect 12716 9911 12768 9920
rect 12716 9877 12725 9911
rect 12725 9877 12759 9911
rect 12759 9877 12768 9911
rect 12716 9868 12768 9877
rect 14188 9868 14240 9920
rect 15844 10004 15896 10056
rect 15936 10004 15988 10056
rect 16856 10047 16908 10056
rect 16856 10013 16865 10047
rect 16865 10013 16899 10047
rect 16899 10013 16908 10047
rect 16856 10004 16908 10013
rect 15660 9868 15712 9920
rect 20812 9936 20864 9988
rect 22008 9936 22060 9988
rect 19892 9911 19944 9920
rect 19892 9877 19901 9911
rect 19901 9877 19935 9911
rect 19935 9877 19944 9911
rect 19892 9868 19944 9877
rect 21272 9911 21324 9920
rect 21272 9877 21281 9911
rect 21281 9877 21315 9911
rect 21315 9877 21324 9911
rect 21272 9868 21324 9877
rect 21364 9868 21416 9920
rect 21916 9911 21968 9920
rect 21916 9877 21925 9911
rect 21925 9877 21959 9911
rect 21959 9877 21968 9911
rect 21916 9868 21968 9877
rect 22560 9868 22612 9920
rect 3662 9766 3714 9818
rect 3726 9766 3778 9818
rect 3790 9766 3842 9818
rect 3854 9766 3906 9818
rect 3918 9766 3970 9818
rect 4620 9707 4672 9716
rect 4620 9673 4629 9707
rect 4629 9673 4663 9707
rect 4663 9673 4672 9707
rect 4620 9664 4672 9673
rect 4988 9596 5040 9648
rect 5080 9596 5132 9648
rect 12716 9664 12768 9716
rect 4712 9571 4764 9580
rect 4712 9537 4721 9571
rect 4721 9537 4755 9571
rect 4755 9537 4764 9571
rect 4712 9528 4764 9537
rect 4804 9528 4856 9580
rect 4896 9503 4948 9512
rect 4896 9469 4905 9503
rect 4905 9469 4939 9503
rect 4939 9469 4948 9503
rect 4896 9460 4948 9469
rect 5448 9503 5500 9512
rect 5448 9469 5457 9503
rect 5457 9469 5491 9503
rect 5491 9469 5500 9503
rect 5448 9460 5500 9469
rect 8852 9571 8904 9580
rect 8852 9537 8861 9571
rect 8861 9537 8895 9571
rect 8895 9537 8904 9571
rect 8852 9528 8904 9537
rect 10508 9571 10560 9580
rect 10508 9537 10517 9571
rect 10517 9537 10551 9571
rect 10551 9537 10560 9571
rect 10508 9528 10560 9537
rect 10692 9571 10744 9580
rect 10692 9537 10701 9571
rect 10701 9537 10735 9571
rect 10735 9537 10744 9571
rect 10692 9528 10744 9537
rect 13912 9664 13964 9716
rect 17408 9707 17460 9716
rect 17408 9673 17417 9707
rect 17417 9673 17451 9707
rect 17451 9673 17460 9707
rect 17408 9664 17460 9673
rect 16856 9596 16908 9648
rect 20812 9707 20864 9716
rect 20812 9673 20821 9707
rect 20821 9673 20855 9707
rect 20855 9673 20864 9707
rect 20812 9664 20864 9673
rect 21364 9664 21416 9716
rect 22468 9664 22520 9716
rect 4712 9392 4764 9444
rect 12900 9503 12952 9512
rect 12900 9469 12909 9503
rect 12909 9469 12943 9503
rect 12943 9469 12952 9503
rect 12900 9460 12952 9469
rect 15384 9528 15436 9580
rect 5724 9324 5776 9376
rect 6276 9324 6328 9376
rect 8392 9367 8444 9376
rect 8392 9333 8401 9367
rect 8401 9333 8435 9367
rect 8435 9333 8444 9367
rect 8392 9324 8444 9333
rect 8760 9367 8812 9376
rect 8760 9333 8769 9367
rect 8769 9333 8803 9367
rect 8803 9333 8812 9367
rect 8760 9324 8812 9333
rect 10048 9367 10100 9376
rect 10048 9333 10057 9367
rect 10057 9333 10091 9367
rect 10091 9333 10100 9367
rect 10048 9324 10100 9333
rect 10784 9324 10836 9376
rect 13636 9460 13688 9512
rect 13820 9503 13872 9512
rect 13820 9469 13854 9503
rect 13854 9469 13872 9503
rect 13820 9460 13872 9469
rect 15752 9460 15804 9512
rect 15844 9503 15896 9512
rect 15844 9469 15853 9503
rect 15853 9469 15887 9503
rect 15887 9469 15896 9503
rect 15844 9460 15896 9469
rect 16488 9460 16540 9512
rect 16580 9503 16632 9512
rect 16580 9469 16589 9503
rect 16589 9469 16623 9503
rect 16623 9469 16632 9503
rect 16580 9460 16632 9469
rect 16672 9503 16724 9512
rect 16672 9469 16681 9503
rect 16681 9469 16715 9503
rect 16715 9469 16724 9503
rect 16672 9460 16724 9469
rect 18144 9528 18196 9580
rect 18052 9460 18104 9512
rect 14096 9324 14148 9376
rect 15660 9367 15712 9376
rect 15660 9333 15669 9367
rect 15669 9333 15703 9367
rect 15703 9333 15712 9367
rect 15660 9324 15712 9333
rect 16856 9324 16908 9376
rect 17500 9324 17552 9376
rect 20904 9503 20956 9512
rect 20904 9469 20913 9503
rect 20913 9469 20947 9503
rect 20947 9469 20956 9503
rect 20904 9460 20956 9469
rect 20720 9392 20772 9444
rect 21180 9528 21232 9580
rect 19156 9367 19208 9376
rect 19156 9333 19165 9367
rect 19165 9333 19199 9367
rect 19199 9333 19208 9367
rect 19156 9324 19208 9333
rect 21272 9392 21324 9444
rect 22468 9324 22520 9376
rect 4322 9222 4374 9274
rect 4386 9222 4438 9274
rect 4450 9222 4502 9274
rect 4514 9222 4566 9274
rect 4578 9222 4630 9274
rect 8760 9120 8812 9172
rect 10784 9163 10836 9172
rect 10784 9129 10793 9163
rect 10793 9129 10827 9163
rect 10827 9129 10836 9163
rect 10784 9120 10836 9129
rect 15660 9120 15712 9172
rect 17408 9120 17460 9172
rect 18144 9163 18196 9172
rect 18144 9129 18153 9163
rect 18153 9129 18187 9163
rect 18187 9129 18196 9163
rect 18144 9120 18196 9129
rect 19340 9120 19392 9172
rect 22560 9120 22612 9172
rect 8392 9052 8444 9104
rect 10048 9052 10100 9104
rect 3056 9027 3108 9036
rect 3056 8993 3065 9027
rect 3065 8993 3099 9027
rect 3099 8993 3108 9027
rect 3056 8984 3108 8993
rect 3332 9027 3384 9036
rect 3332 8993 3341 9027
rect 3341 8993 3375 9027
rect 3375 8993 3384 9027
rect 3332 8984 3384 8993
rect 3516 8916 3568 8968
rect 4160 8984 4212 9036
rect 4988 8984 5040 9036
rect 8852 8984 8904 9036
rect 9404 9027 9456 9036
rect 9404 8993 9413 9027
rect 9413 8993 9447 9027
rect 9447 8993 9456 9027
rect 9404 8984 9456 8993
rect 11428 9027 11480 9036
rect 11428 8993 11437 9027
rect 11437 8993 11471 9027
rect 11471 8993 11480 9027
rect 11428 8984 11480 8993
rect 12900 9052 12952 9104
rect 14096 9027 14148 9036
rect 14096 8993 14105 9027
rect 14105 8993 14139 9027
rect 14139 8993 14148 9027
rect 14096 8984 14148 8993
rect 19156 9052 19208 9104
rect 15568 9027 15620 9036
rect 15568 8993 15577 9027
rect 15577 8993 15611 9027
rect 15611 8993 15620 9027
rect 15568 8984 15620 8993
rect 4068 8959 4120 8968
rect 4068 8925 4077 8959
rect 4077 8925 4111 8959
rect 4111 8925 4120 8959
rect 4068 8916 4120 8925
rect 11244 8916 11296 8968
rect 11612 8916 11664 8968
rect 13912 8916 13964 8968
rect 13820 8848 13872 8900
rect 14004 8848 14056 8900
rect 15752 8848 15804 8900
rect 17500 9027 17552 9036
rect 17500 8993 17518 9027
rect 17518 8993 17552 9027
rect 17500 8984 17552 8993
rect 21364 8984 21416 9036
rect 16672 8848 16724 8900
rect 3148 8823 3200 8832
rect 3148 8789 3157 8823
rect 3157 8789 3191 8823
rect 3191 8789 3200 8823
rect 3148 8780 3200 8789
rect 4068 8780 4120 8832
rect 5080 8823 5132 8832
rect 5080 8789 5089 8823
rect 5089 8789 5123 8823
rect 5123 8789 5132 8823
rect 5080 8780 5132 8789
rect 5908 8780 5960 8832
rect 10968 8780 11020 8832
rect 12532 8780 12584 8832
rect 14188 8823 14240 8832
rect 14188 8789 14197 8823
rect 14197 8789 14231 8823
rect 14231 8789 14240 8823
rect 14188 8780 14240 8789
rect 20812 8916 20864 8968
rect 20812 8780 20864 8832
rect 3662 8678 3714 8730
rect 3726 8678 3778 8730
rect 3790 8678 3842 8730
rect 3854 8678 3906 8730
rect 3918 8678 3970 8730
rect 4068 8576 4120 8628
rect 4988 8619 5040 8628
rect 4988 8585 4997 8619
rect 4997 8585 5031 8619
rect 5031 8585 5040 8619
rect 4988 8576 5040 8585
rect 5724 8576 5776 8628
rect 6368 8576 6420 8628
rect 5448 8508 5500 8560
rect 6092 8508 6144 8560
rect 3148 8372 3200 8424
rect 3424 8304 3476 8356
rect 6276 8415 6328 8424
rect 6276 8381 6285 8415
rect 6285 8381 6319 8415
rect 6319 8381 6328 8415
rect 6276 8372 6328 8381
rect 6368 8415 6420 8424
rect 6368 8381 6377 8415
rect 6377 8381 6411 8415
rect 6411 8381 6420 8415
rect 6368 8372 6420 8381
rect 6736 8372 6788 8424
rect 7748 8619 7800 8628
rect 7748 8585 7757 8619
rect 7757 8585 7791 8619
rect 7791 8585 7800 8619
rect 7748 8576 7800 8585
rect 10968 8576 11020 8628
rect 15476 8619 15528 8628
rect 15476 8585 15485 8619
rect 15485 8585 15519 8619
rect 15519 8585 15528 8619
rect 15476 8576 15528 8585
rect 16672 8576 16724 8628
rect 21364 8576 21416 8628
rect 22008 8576 22060 8628
rect 11152 8508 11204 8560
rect 4160 8304 4212 8356
rect 4712 8304 4764 8356
rect 4804 8347 4856 8356
rect 4804 8313 4829 8347
rect 4829 8313 4856 8347
rect 4804 8304 4856 8313
rect 5816 8347 5868 8356
rect 5816 8313 5825 8347
rect 5825 8313 5859 8347
rect 5859 8313 5868 8347
rect 5816 8304 5868 8313
rect 6184 8279 6236 8288
rect 6184 8245 6193 8279
rect 6193 8245 6227 8279
rect 6227 8245 6236 8279
rect 6184 8236 6236 8245
rect 7748 8236 7800 8288
rect 8208 8236 8260 8288
rect 8760 8440 8812 8492
rect 10784 8440 10836 8492
rect 11428 8415 11480 8424
rect 11428 8381 11437 8415
rect 11437 8381 11471 8415
rect 11471 8381 11480 8415
rect 11428 8372 11480 8381
rect 11612 8415 11664 8424
rect 11612 8381 11621 8415
rect 11621 8381 11655 8415
rect 11655 8381 11664 8415
rect 11612 8372 11664 8381
rect 12532 8415 12584 8424
rect 12532 8381 12541 8415
rect 12541 8381 12575 8415
rect 12575 8381 12584 8415
rect 12532 8372 12584 8381
rect 12900 8372 12952 8424
rect 13544 8440 13596 8492
rect 14188 8440 14240 8492
rect 21916 8508 21968 8560
rect 14096 8372 14148 8424
rect 14188 8347 14240 8356
rect 14188 8313 14197 8347
rect 14197 8313 14231 8347
rect 14231 8313 14240 8347
rect 14188 8304 14240 8313
rect 15752 8415 15804 8424
rect 15752 8381 15761 8415
rect 15761 8381 15795 8415
rect 15795 8381 15804 8415
rect 15752 8372 15804 8381
rect 15568 8304 15620 8356
rect 16212 8304 16264 8356
rect 20996 8304 21048 8356
rect 21272 8304 21324 8356
rect 11612 8236 11664 8288
rect 12808 8236 12860 8288
rect 14464 8236 14516 8288
rect 15384 8236 15436 8288
rect 19156 8236 19208 8288
rect 4322 8134 4374 8186
rect 4386 8134 4438 8186
rect 4450 8134 4502 8186
rect 4514 8134 4566 8186
rect 4578 8134 4630 8186
rect 3148 8032 3200 8084
rect 3516 8032 3568 8084
rect 4712 8032 4764 8084
rect 3056 7964 3108 8016
rect 15476 8032 15528 8084
rect 16212 8032 16264 8084
rect 16856 8075 16908 8084
rect 16856 8041 16883 8075
rect 16883 8041 16908 8075
rect 16856 8032 16908 8041
rect 21456 8032 21508 8084
rect 3148 7939 3200 7948
rect 3148 7905 3157 7939
rect 3157 7905 3191 7939
rect 3191 7905 3200 7939
rect 3148 7896 3200 7905
rect 3332 7939 3384 7948
rect 3332 7905 3341 7939
rect 3341 7905 3375 7939
rect 3375 7905 3384 7939
rect 3332 7896 3384 7905
rect 3424 7939 3476 7948
rect 3424 7905 3433 7939
rect 3433 7905 3467 7939
rect 3467 7905 3476 7939
rect 3424 7896 3476 7905
rect 5908 7939 5960 7948
rect 5908 7905 5917 7939
rect 5917 7905 5951 7939
rect 5951 7905 5960 7939
rect 5908 7896 5960 7905
rect 6184 7896 6236 7948
rect 6736 7896 6788 7948
rect 8392 7896 8444 7948
rect 8760 7896 8812 7948
rect 10968 7896 11020 7948
rect 11612 7939 11664 7948
rect 11612 7905 11621 7939
rect 11621 7905 11655 7939
rect 11655 7905 11664 7939
rect 11612 7896 11664 7905
rect 6368 7828 6420 7880
rect 7380 7828 7432 7880
rect 8208 7828 8260 7880
rect 11152 7828 11204 7880
rect 13544 7939 13596 7948
rect 13544 7905 13553 7939
rect 13553 7905 13587 7939
rect 13587 7905 13596 7939
rect 13544 7896 13596 7905
rect 14188 7964 14240 8016
rect 16488 8007 16540 8016
rect 16488 7973 16497 8007
rect 16497 7973 16531 8007
rect 16531 7973 16540 8007
rect 16488 7964 16540 7973
rect 13912 7896 13964 7948
rect 14280 7939 14332 7948
rect 14280 7905 14289 7939
rect 14289 7905 14323 7939
rect 14323 7905 14332 7939
rect 14280 7896 14332 7905
rect 13268 7828 13320 7880
rect 16856 7896 16908 7948
rect 18328 7896 18380 7948
rect 19248 7964 19300 8016
rect 18788 7896 18840 7948
rect 21824 7964 21876 8016
rect 21916 7939 21968 7948
rect 21916 7905 21925 7939
rect 21925 7905 21959 7939
rect 21959 7905 21968 7939
rect 21916 7896 21968 7905
rect 16672 7828 16724 7880
rect 21456 7871 21508 7880
rect 21456 7837 21465 7871
rect 21465 7837 21499 7871
rect 21499 7837 21508 7871
rect 21456 7828 21508 7837
rect 9496 7760 9548 7812
rect 2320 7735 2372 7744
rect 2320 7701 2329 7735
rect 2329 7701 2363 7735
rect 2363 7701 2372 7735
rect 2320 7692 2372 7701
rect 2412 7692 2464 7744
rect 2964 7735 3016 7744
rect 2964 7701 2973 7735
rect 2973 7701 3007 7735
rect 3007 7701 3016 7735
rect 2964 7692 3016 7701
rect 4252 7692 4304 7744
rect 6092 7735 6144 7744
rect 6092 7701 6101 7735
rect 6101 7701 6135 7735
rect 6135 7701 6144 7735
rect 6092 7692 6144 7701
rect 6920 7735 6972 7744
rect 6920 7701 6929 7735
rect 6929 7701 6963 7735
rect 6963 7701 6972 7735
rect 6920 7692 6972 7701
rect 7932 7735 7984 7744
rect 7932 7701 7941 7735
rect 7941 7701 7975 7735
rect 7975 7701 7984 7735
rect 7932 7692 7984 7701
rect 9772 7692 9824 7744
rect 11060 7735 11112 7744
rect 11060 7701 11069 7735
rect 11069 7701 11103 7735
rect 11103 7701 11112 7735
rect 11060 7692 11112 7701
rect 11612 7735 11664 7744
rect 11612 7701 11621 7735
rect 11621 7701 11655 7735
rect 11655 7701 11664 7735
rect 11612 7692 11664 7701
rect 13636 7692 13688 7744
rect 14004 7735 14056 7744
rect 14004 7701 14013 7735
rect 14013 7701 14047 7735
rect 14047 7701 14056 7735
rect 14004 7692 14056 7701
rect 16580 7692 16632 7744
rect 19892 7760 19944 7812
rect 22836 7828 22888 7880
rect 21364 7692 21416 7744
rect 3662 7590 3714 7642
rect 3726 7590 3778 7642
rect 3790 7590 3842 7642
rect 3854 7590 3906 7642
rect 3918 7590 3970 7642
rect 3148 7488 3200 7540
rect 7380 7531 7432 7540
rect 7380 7497 7389 7531
rect 7389 7497 7423 7531
rect 7423 7497 7432 7531
rect 7380 7488 7432 7497
rect 7932 7531 7984 7540
rect 7932 7497 7941 7531
rect 7941 7497 7975 7531
rect 7975 7497 7984 7531
rect 7932 7488 7984 7497
rect 8392 7531 8444 7540
rect 8392 7497 8401 7531
rect 8401 7497 8435 7531
rect 8435 7497 8444 7531
rect 8392 7488 8444 7497
rect 8208 7420 8260 7472
rect 13268 7531 13320 7540
rect 13268 7497 13277 7531
rect 13277 7497 13311 7531
rect 13311 7497 13320 7531
rect 13268 7488 13320 7497
rect 14004 7531 14056 7540
rect 14004 7497 14013 7531
rect 14013 7497 14047 7531
rect 14047 7497 14056 7531
rect 14004 7488 14056 7497
rect 14280 7531 14332 7540
rect 14280 7497 14289 7531
rect 14289 7497 14323 7531
rect 14323 7497 14332 7531
rect 14280 7488 14332 7497
rect 18788 7531 18840 7540
rect 18788 7497 18797 7531
rect 18797 7497 18831 7531
rect 18831 7497 18840 7531
rect 18788 7488 18840 7497
rect 20720 7531 20772 7540
rect 20720 7497 20729 7531
rect 20729 7497 20763 7531
rect 20763 7497 20772 7531
rect 20720 7488 20772 7497
rect 21364 7531 21416 7540
rect 21364 7497 21373 7531
rect 21373 7497 21407 7531
rect 21407 7497 21416 7531
rect 21364 7488 21416 7497
rect 2872 7352 2924 7404
rect 3240 7395 3292 7404
rect 3240 7361 3249 7395
rect 3249 7361 3283 7395
rect 3283 7361 3292 7395
rect 3240 7352 3292 7361
rect 4712 7352 4764 7404
rect 6920 7352 6972 7404
rect 3056 7284 3108 7336
rect 4896 7327 4948 7336
rect 4896 7293 4905 7327
rect 4905 7293 4939 7327
rect 4939 7293 4948 7327
rect 4896 7284 4948 7293
rect 7196 7284 7248 7336
rect 11612 7352 11664 7404
rect 12808 7395 12860 7404
rect 12808 7361 12817 7395
rect 12817 7361 12851 7395
rect 12851 7361 12860 7395
rect 12808 7352 12860 7361
rect 13636 7395 13688 7404
rect 13636 7361 13645 7395
rect 13645 7361 13679 7395
rect 13679 7361 13688 7395
rect 13636 7352 13688 7361
rect 14464 7395 14516 7404
rect 14464 7361 14473 7395
rect 14473 7361 14507 7395
rect 14507 7361 14516 7395
rect 14464 7352 14516 7361
rect 8208 7327 8260 7336
rect 8208 7293 8217 7327
rect 8217 7293 8251 7327
rect 8251 7293 8260 7327
rect 8208 7284 8260 7293
rect 10692 7327 10744 7336
rect 10692 7293 10701 7327
rect 10701 7293 10735 7327
rect 10735 7293 10744 7327
rect 10692 7284 10744 7293
rect 12992 7284 13044 7336
rect 13820 7284 13872 7336
rect 14556 7327 14608 7336
rect 14556 7293 14565 7327
rect 14565 7293 14599 7327
rect 14599 7293 14608 7327
rect 14556 7284 14608 7293
rect 15568 7284 15620 7336
rect 16856 7352 16908 7404
rect 16488 7284 16540 7336
rect 19432 7352 19484 7404
rect 2136 7216 2188 7268
rect 3700 7216 3752 7268
rect 7656 7216 7708 7268
rect 19156 7259 19208 7268
rect 19156 7225 19165 7259
rect 19165 7225 19199 7259
rect 19199 7225 19208 7259
rect 19156 7216 19208 7225
rect 19892 7352 19944 7404
rect 19800 7284 19852 7336
rect 19984 7216 20036 7268
rect 21916 7352 21968 7404
rect 22192 7395 22244 7404
rect 22192 7361 22201 7395
rect 22201 7361 22235 7395
rect 22235 7361 22244 7395
rect 22192 7352 22244 7361
rect 22376 7352 22428 7404
rect 20996 7327 21048 7336
rect 20996 7293 21005 7327
rect 21005 7293 21039 7327
rect 21039 7293 21048 7327
rect 20996 7284 21048 7293
rect 22468 7327 22520 7336
rect 22468 7293 22477 7327
rect 22477 7293 22511 7327
rect 22511 7293 22520 7327
rect 22468 7284 22520 7293
rect 21824 7216 21876 7268
rect 3332 7148 3384 7200
rect 3608 7148 3660 7200
rect 4804 7148 4856 7200
rect 8208 7148 8260 7200
rect 11612 7148 11664 7200
rect 16212 7191 16264 7200
rect 16212 7157 16221 7191
rect 16221 7157 16255 7191
rect 16255 7157 16264 7191
rect 16212 7148 16264 7157
rect 19340 7148 19392 7200
rect 20536 7191 20588 7200
rect 20536 7157 20545 7191
rect 20545 7157 20579 7191
rect 20579 7157 20588 7191
rect 20536 7148 20588 7157
rect 21272 7148 21324 7200
rect 21548 7191 21600 7200
rect 21548 7157 21557 7191
rect 21557 7157 21591 7191
rect 21591 7157 21600 7191
rect 21548 7148 21600 7157
rect 4322 7046 4374 7098
rect 4386 7046 4438 7098
rect 4450 7046 4502 7098
rect 4514 7046 4566 7098
rect 4578 7046 4630 7098
rect 2136 6987 2188 6996
rect 2136 6953 2145 6987
rect 2145 6953 2179 6987
rect 2179 6953 2188 6987
rect 2136 6944 2188 6953
rect 2412 6944 2464 6996
rect 3056 6944 3108 6996
rect 2780 6876 2832 6928
rect 3700 6944 3752 6996
rect 4896 6944 4948 6996
rect 3424 6919 3476 6928
rect 3424 6885 3451 6919
rect 3451 6885 3476 6919
rect 3424 6876 3476 6885
rect 3608 6919 3660 6928
rect 3608 6885 3617 6919
rect 3617 6885 3651 6919
rect 3651 6885 3660 6919
rect 3608 6876 3660 6885
rect 9772 6876 9824 6928
rect 4804 6808 4856 6860
rect 10048 6808 10100 6860
rect 11152 6851 11204 6860
rect 11152 6817 11161 6851
rect 11161 6817 11195 6851
rect 11195 6817 11204 6851
rect 11152 6808 11204 6817
rect 15568 6919 15620 6928
rect 15568 6885 15577 6919
rect 15577 6885 15611 6919
rect 15611 6885 15620 6919
rect 15568 6876 15620 6885
rect 16488 6876 16540 6928
rect 21456 6944 21508 6996
rect 19984 6876 20036 6928
rect 16396 6851 16448 6860
rect 16396 6817 16430 6851
rect 16430 6817 16448 6851
rect 5632 6783 5684 6792
rect 5632 6749 5641 6783
rect 5641 6749 5675 6783
rect 5675 6749 5684 6783
rect 5632 6740 5684 6749
rect 9496 6783 9548 6792
rect 9496 6749 9505 6783
rect 9505 6749 9539 6783
rect 9539 6749 9548 6783
rect 9496 6740 9548 6749
rect 11060 6783 11112 6792
rect 11060 6749 11069 6783
rect 11069 6749 11103 6783
rect 11103 6749 11112 6783
rect 11060 6740 11112 6749
rect 16396 6808 16448 6817
rect 18328 6851 18380 6860
rect 18328 6817 18337 6851
rect 18337 6817 18371 6851
rect 18371 6817 18380 6851
rect 18328 6808 18380 6817
rect 18604 6851 18656 6860
rect 18604 6817 18638 6851
rect 18638 6817 18656 6851
rect 18604 6808 18656 6817
rect 19892 6851 19944 6860
rect 19892 6817 19901 6851
rect 19901 6817 19935 6851
rect 19935 6817 19944 6851
rect 19892 6808 19944 6817
rect 21548 6876 21600 6928
rect 15936 6740 15988 6792
rect 13912 6672 13964 6724
rect 19708 6715 19760 6724
rect 19708 6681 19717 6715
rect 19717 6681 19751 6715
rect 19751 6681 19760 6715
rect 20260 6808 20312 6860
rect 21180 6808 21232 6860
rect 19708 6672 19760 6681
rect 2320 6647 2372 6656
rect 2320 6613 2329 6647
rect 2329 6613 2363 6647
rect 2363 6613 2372 6647
rect 2320 6604 2372 6613
rect 2964 6647 3016 6656
rect 2964 6613 2973 6647
rect 2973 6613 3007 6647
rect 3007 6613 3016 6647
rect 2964 6604 3016 6613
rect 3240 6604 3292 6656
rect 11612 6647 11664 6656
rect 11612 6613 11621 6647
rect 11621 6613 11655 6647
rect 11655 6613 11664 6647
rect 11612 6604 11664 6613
rect 16120 6604 16172 6656
rect 19984 6604 20036 6656
rect 20904 6740 20956 6792
rect 21272 6740 21324 6792
rect 20720 6672 20772 6724
rect 21272 6604 21324 6656
rect 21824 6604 21876 6656
rect 3662 6502 3714 6554
rect 3726 6502 3778 6554
rect 3790 6502 3842 6554
rect 3854 6502 3906 6554
rect 3918 6502 3970 6554
rect 4712 6400 4764 6452
rect 4804 6443 4856 6452
rect 4804 6409 4813 6443
rect 4813 6409 4847 6443
rect 4847 6409 4856 6443
rect 4804 6400 4856 6409
rect 13820 6443 13872 6452
rect 13820 6409 13829 6443
rect 13829 6409 13863 6443
rect 13863 6409 13872 6443
rect 13820 6400 13872 6409
rect 14280 6400 14332 6452
rect 15568 6400 15620 6452
rect 16212 6443 16264 6452
rect 16212 6409 16221 6443
rect 16221 6409 16255 6443
rect 16255 6409 16264 6443
rect 16212 6400 16264 6409
rect 16396 6443 16448 6452
rect 16396 6409 16405 6443
rect 16405 6409 16439 6443
rect 16439 6409 16448 6443
rect 16396 6400 16448 6409
rect 18604 6400 18656 6452
rect 19156 6400 19208 6452
rect 19432 6400 19484 6452
rect 19800 6443 19852 6452
rect 19800 6409 19809 6443
rect 19809 6409 19843 6443
rect 19843 6409 19852 6443
rect 19800 6400 19852 6409
rect 19984 6443 20036 6452
rect 19984 6409 19993 6443
rect 19993 6409 20027 6443
rect 20027 6409 20036 6443
rect 19984 6400 20036 6409
rect 20904 6400 20956 6452
rect 4252 6375 4304 6384
rect 4252 6341 4261 6375
rect 4261 6341 4295 6375
rect 4295 6341 4304 6375
rect 4252 6332 4304 6341
rect 5816 6332 5868 6384
rect 6828 6332 6880 6384
rect 5816 6196 5868 6248
rect 6736 6264 6788 6316
rect 6552 6196 6604 6248
rect 3516 6060 3568 6112
rect 7196 6196 7248 6248
rect 11980 6332 12032 6384
rect 22100 6400 22152 6452
rect 19432 6264 19484 6316
rect 19708 6307 19760 6316
rect 19708 6273 19717 6307
rect 19717 6273 19751 6307
rect 19751 6273 19760 6307
rect 19708 6264 19760 6273
rect 20536 6264 20588 6316
rect 7380 6239 7432 6248
rect 7380 6205 7389 6239
rect 7389 6205 7423 6239
rect 7423 6205 7432 6239
rect 7380 6196 7432 6205
rect 7656 6239 7708 6248
rect 7656 6205 7665 6239
rect 7665 6205 7699 6239
rect 7699 6205 7708 6239
rect 7656 6196 7708 6205
rect 14556 6196 14608 6248
rect 19340 6196 19392 6248
rect 19800 6196 19852 6248
rect 12992 6128 13044 6180
rect 13728 6128 13780 6180
rect 5540 6103 5592 6112
rect 5540 6069 5549 6103
rect 5549 6069 5583 6103
rect 5583 6069 5592 6103
rect 5540 6060 5592 6069
rect 5724 6103 5776 6112
rect 5724 6069 5751 6103
rect 5751 6069 5776 6103
rect 5724 6060 5776 6069
rect 6368 6060 6420 6112
rect 6460 6103 6512 6112
rect 6460 6069 6469 6103
rect 6469 6069 6503 6103
rect 6503 6069 6512 6103
rect 6460 6060 6512 6069
rect 6736 6060 6788 6112
rect 7380 6060 7432 6112
rect 8024 6060 8076 6112
rect 13360 6060 13412 6112
rect 14004 6103 14056 6112
rect 14004 6069 14013 6103
rect 14013 6069 14047 6103
rect 14047 6069 14056 6103
rect 14924 6171 14976 6180
rect 14924 6137 14933 6171
rect 14933 6137 14967 6171
rect 14967 6137 14976 6171
rect 14924 6128 14976 6137
rect 16028 6171 16080 6180
rect 16028 6137 16037 6171
rect 16037 6137 16071 6171
rect 16071 6137 16080 6171
rect 16028 6128 16080 6137
rect 16120 6128 16172 6180
rect 21088 6196 21140 6248
rect 20260 6128 20312 6180
rect 14004 6060 14056 6069
rect 14280 6103 14332 6112
rect 14280 6069 14289 6103
rect 14289 6069 14323 6103
rect 14323 6069 14332 6103
rect 14280 6060 14332 6069
rect 14556 6060 14608 6112
rect 15200 6060 15252 6112
rect 15936 6060 15988 6112
rect 16488 6060 16540 6112
rect 20812 6128 20864 6180
rect 22560 6196 22612 6248
rect 22836 6103 22888 6112
rect 22836 6069 22845 6103
rect 22845 6069 22879 6103
rect 22879 6069 22888 6103
rect 22836 6060 22888 6069
rect 4322 5958 4374 6010
rect 4386 5958 4438 6010
rect 4450 5958 4502 6010
rect 4514 5958 4566 6010
rect 4578 5958 4630 6010
rect 5724 5856 5776 5908
rect 7196 5856 7248 5908
rect 7656 5856 7708 5908
rect 4252 5788 4304 5840
rect 5816 5788 5868 5840
rect 6736 5788 6788 5840
rect 6368 5763 6420 5772
rect 6368 5729 6402 5763
rect 6402 5729 6420 5763
rect 6368 5720 6420 5729
rect 8300 5720 8352 5772
rect 8852 5720 8904 5772
rect 9404 5856 9456 5908
rect 10048 5788 10100 5840
rect 5632 5652 5684 5704
rect 9864 5763 9916 5772
rect 9864 5729 9873 5763
rect 9873 5729 9907 5763
rect 9907 5729 9916 5763
rect 9864 5720 9916 5729
rect 10232 5831 10284 5840
rect 10232 5797 10241 5831
rect 10241 5797 10275 5831
rect 10275 5797 10284 5831
rect 10232 5788 10284 5797
rect 11152 5856 11204 5908
rect 11980 5899 12032 5908
rect 11980 5865 11989 5899
rect 11989 5865 12023 5899
rect 12023 5865 12032 5899
rect 11980 5856 12032 5865
rect 13728 5856 13780 5908
rect 19984 5899 20036 5908
rect 19984 5865 19993 5899
rect 19993 5865 20027 5899
rect 20027 5865 20036 5899
rect 19984 5856 20036 5865
rect 20260 5856 20312 5908
rect 20996 5856 21048 5908
rect 12532 5788 12584 5840
rect 15384 5788 15436 5840
rect 16028 5788 16080 5840
rect 10692 5720 10744 5772
rect 12992 5763 13044 5772
rect 12992 5729 13001 5763
rect 13001 5729 13035 5763
rect 13035 5729 13044 5763
rect 12992 5720 13044 5729
rect 11428 5652 11480 5704
rect 14004 5763 14056 5772
rect 14004 5729 14013 5763
rect 14013 5729 14047 5763
rect 14047 5729 14056 5763
rect 14004 5720 14056 5729
rect 14280 5763 14332 5772
rect 14280 5729 14289 5763
rect 14289 5729 14323 5763
rect 14323 5729 14332 5763
rect 14280 5720 14332 5729
rect 14556 5763 14608 5772
rect 14556 5729 14565 5763
rect 14565 5729 14599 5763
rect 14599 5729 14608 5763
rect 14556 5720 14608 5729
rect 15568 5720 15620 5772
rect 18328 5720 18380 5772
rect 19708 5788 19760 5840
rect 18880 5763 18932 5772
rect 18880 5729 18914 5763
rect 18914 5729 18932 5763
rect 18880 5720 18932 5729
rect 22560 5899 22612 5908
rect 22560 5865 22569 5899
rect 22569 5865 22603 5899
rect 22603 5865 22612 5899
rect 22560 5856 22612 5865
rect 20352 5720 20404 5772
rect 20628 5720 20680 5772
rect 21272 5763 21324 5772
rect 21272 5729 21281 5763
rect 21281 5729 21315 5763
rect 21315 5729 21324 5763
rect 21272 5720 21324 5729
rect 21824 5720 21876 5772
rect 21916 5763 21968 5772
rect 21916 5729 21925 5763
rect 21925 5729 21959 5763
rect 21959 5729 21968 5763
rect 21916 5720 21968 5729
rect 13360 5652 13412 5704
rect 20720 5652 20772 5704
rect 22836 5720 22888 5772
rect 13820 5584 13872 5636
rect 8760 5516 8812 5568
rect 10324 5516 10376 5568
rect 11980 5559 12032 5568
rect 11980 5525 11989 5559
rect 11989 5525 12023 5559
rect 12023 5525 12032 5559
rect 11980 5516 12032 5525
rect 12072 5516 12124 5568
rect 12716 5516 12768 5568
rect 15200 5559 15252 5568
rect 15200 5525 15209 5559
rect 15209 5525 15243 5559
rect 15243 5525 15252 5559
rect 15200 5516 15252 5525
rect 15384 5559 15436 5568
rect 15384 5525 15393 5559
rect 15393 5525 15427 5559
rect 15427 5525 15436 5559
rect 15384 5516 15436 5525
rect 20076 5559 20128 5568
rect 20076 5525 20085 5559
rect 20085 5525 20119 5559
rect 20119 5525 20128 5559
rect 20076 5516 20128 5525
rect 22284 5584 22336 5636
rect 3662 5414 3714 5466
rect 3726 5414 3778 5466
rect 3790 5414 3842 5466
rect 3854 5414 3906 5466
rect 3918 5414 3970 5466
rect 2780 5312 2832 5364
rect 3516 5355 3568 5364
rect 3516 5321 3525 5355
rect 3525 5321 3559 5355
rect 3559 5321 3568 5355
rect 3516 5312 3568 5321
rect 3424 5244 3476 5296
rect 3884 5244 3936 5296
rect 2872 5108 2924 5160
rect 5632 5312 5684 5364
rect 6828 5355 6880 5364
rect 6828 5321 6837 5355
rect 6837 5321 6871 5355
rect 6871 5321 6880 5355
rect 6828 5312 6880 5321
rect 8024 5355 8076 5364
rect 8024 5321 8033 5355
rect 8033 5321 8067 5355
rect 8067 5321 8076 5355
rect 8024 5312 8076 5321
rect 8300 5312 8352 5364
rect 8760 5355 8812 5364
rect 8760 5321 8769 5355
rect 8769 5321 8803 5355
rect 8803 5321 8812 5355
rect 8760 5312 8812 5321
rect 10692 5312 10744 5364
rect 11152 5312 11204 5364
rect 12716 5355 12768 5364
rect 12716 5321 12725 5355
rect 12725 5321 12759 5355
rect 12759 5321 12768 5355
rect 12716 5312 12768 5321
rect 14924 5312 14976 5364
rect 18880 5312 18932 5364
rect 19156 5312 19208 5364
rect 20812 5312 20864 5364
rect 5540 5108 5592 5160
rect 7196 5151 7248 5160
rect 7196 5117 7205 5151
rect 7205 5117 7239 5151
rect 7239 5117 7248 5151
rect 7196 5108 7248 5117
rect 7564 5108 7616 5160
rect 8852 5176 8904 5228
rect 12992 5176 13044 5228
rect 9404 5151 9456 5160
rect 9404 5117 9413 5151
rect 9413 5117 9447 5151
rect 9447 5117 9456 5151
rect 9404 5108 9456 5117
rect 12072 5151 12124 5160
rect 12072 5117 12090 5151
rect 12090 5117 12124 5151
rect 12072 5108 12124 5117
rect 3332 5083 3384 5092
rect 3332 5049 3341 5083
rect 3341 5049 3375 5083
rect 3375 5049 3384 5083
rect 3332 5040 3384 5049
rect 6460 5040 6512 5092
rect 8024 5083 8076 5092
rect 8024 5049 8033 5083
rect 8033 5049 8067 5083
rect 8067 5049 8076 5083
rect 8024 5040 8076 5049
rect 8576 5083 8628 5092
rect 8576 5049 8585 5083
rect 8585 5049 8619 5083
rect 8619 5049 8628 5083
rect 8576 5040 8628 5049
rect 2504 5015 2556 5024
rect 2504 4981 2513 5015
rect 2513 4981 2547 5015
rect 2547 4981 2556 5015
rect 2504 4972 2556 4981
rect 3240 4972 3292 5024
rect 3424 4972 3476 5024
rect 3700 5015 3752 5024
rect 3700 4981 3709 5015
rect 3709 4981 3743 5015
rect 3743 4981 3752 5015
rect 3700 4972 3752 4981
rect 7380 5015 7432 5024
rect 7380 4981 7389 5015
rect 7389 4981 7423 5015
rect 7423 4981 7432 5015
rect 7380 4972 7432 4981
rect 8944 5015 8996 5024
rect 8944 4981 8953 5015
rect 8953 4981 8987 5015
rect 8987 4981 8996 5015
rect 8944 4972 8996 4981
rect 10140 5040 10192 5092
rect 11428 5040 11480 5092
rect 12900 5108 12952 5160
rect 16488 5219 16540 5228
rect 16488 5185 16497 5219
rect 16497 5185 16531 5219
rect 16531 5185 16540 5219
rect 16488 5176 16540 5185
rect 19800 5244 19852 5296
rect 12532 5083 12584 5092
rect 12532 5049 12541 5083
rect 12541 5049 12575 5083
rect 12575 5049 12584 5083
rect 12532 5040 12584 5049
rect 13360 5151 13412 5160
rect 13360 5117 13369 5151
rect 13369 5117 13403 5151
rect 13403 5117 13412 5151
rect 13360 5108 13412 5117
rect 13820 5151 13872 5160
rect 13820 5117 13854 5151
rect 13854 5117 13872 5151
rect 13820 5108 13872 5117
rect 15384 5108 15436 5160
rect 20260 5151 20312 5160
rect 20260 5117 20269 5151
rect 20269 5117 20303 5151
rect 20303 5117 20312 5151
rect 20260 5108 20312 5117
rect 20352 5151 20404 5160
rect 20352 5117 20361 5151
rect 20361 5117 20395 5151
rect 20395 5117 20404 5151
rect 20352 5108 20404 5117
rect 20076 5040 20128 5092
rect 10048 4972 10100 5024
rect 12900 5015 12952 5024
rect 12900 4981 12909 5015
rect 12909 4981 12943 5015
rect 12943 4981 12952 5015
rect 12900 4972 12952 4981
rect 14280 4972 14332 5024
rect 19984 5015 20036 5024
rect 19984 4981 19993 5015
rect 19993 4981 20027 5015
rect 20027 4981 20036 5015
rect 19984 4972 20036 4981
rect 20720 5151 20772 5160
rect 20720 5117 20729 5151
rect 20729 5117 20763 5151
rect 20763 5117 20772 5151
rect 20720 5108 20772 5117
rect 20904 5151 20956 5160
rect 20904 5117 20913 5151
rect 20913 5117 20947 5151
rect 20947 5117 20956 5151
rect 20904 5108 20956 5117
rect 22192 5108 22244 5160
rect 4322 4870 4374 4922
rect 4386 4870 4438 4922
rect 4450 4870 4502 4922
rect 4514 4870 4566 4922
rect 4578 4870 4630 4922
rect 4068 4768 4120 4820
rect 6552 4811 6604 4820
rect 6552 4777 6561 4811
rect 6561 4777 6595 4811
rect 6595 4777 6604 4811
rect 6552 4768 6604 4777
rect 8024 4811 8076 4820
rect 8024 4777 8033 4811
rect 8033 4777 8067 4811
rect 8067 4777 8076 4811
rect 8024 4768 8076 4777
rect 2504 4700 2556 4752
rect 2872 4700 2924 4752
rect 3884 4743 3936 4752
rect 3884 4709 3893 4743
rect 3893 4709 3927 4743
rect 3927 4709 3936 4743
rect 3884 4700 3936 4709
rect 4712 4743 4764 4752
rect 4712 4709 4739 4743
rect 4739 4709 4764 4743
rect 4712 4700 4764 4709
rect 5632 4700 5684 4752
rect 5724 4700 5776 4752
rect 1676 4632 1728 4684
rect 3056 4632 3108 4684
rect 3148 4632 3200 4684
rect 4160 4632 4212 4684
rect 2320 4607 2372 4616
rect 2320 4573 2329 4607
rect 2329 4573 2363 4607
rect 2363 4573 2372 4607
rect 2320 4564 2372 4573
rect 1768 4428 1820 4480
rect 2780 4428 2832 4480
rect 4436 4539 4488 4548
rect 4436 4505 4445 4539
rect 4445 4505 4479 4539
rect 4479 4505 4488 4539
rect 4436 4496 4488 4505
rect 4344 4428 4396 4480
rect 6828 4700 6880 4752
rect 8576 4768 8628 4820
rect 8944 4743 8996 4752
rect 8944 4709 8978 4743
rect 8978 4709 8996 4743
rect 8944 4700 8996 4709
rect 10140 4811 10192 4820
rect 10140 4777 10149 4811
rect 10149 4777 10183 4811
rect 10183 4777 10192 4811
rect 10140 4768 10192 4777
rect 11888 4768 11940 4820
rect 13728 4768 13780 4820
rect 20260 4768 20312 4820
rect 20904 4768 20956 4820
rect 12900 4700 12952 4752
rect 19984 4743 20036 4752
rect 19984 4709 20018 4743
rect 20018 4709 20036 4743
rect 19984 4700 20036 4709
rect 7380 4564 7432 4616
rect 8760 4632 8812 4684
rect 11428 4632 11480 4684
rect 12808 4607 12860 4616
rect 12808 4573 12817 4607
rect 12817 4573 12851 4607
rect 12851 4573 12860 4607
rect 12808 4564 12860 4573
rect 19708 4607 19760 4616
rect 19708 4573 19717 4607
rect 19717 4573 19751 4607
rect 19751 4573 19760 4607
rect 19708 4564 19760 4573
rect 10232 4496 10284 4548
rect 7196 4428 7248 4480
rect 10048 4471 10100 4480
rect 10048 4437 10057 4471
rect 10057 4437 10091 4471
rect 10091 4437 10100 4471
rect 10048 4428 10100 4437
rect 10324 4471 10376 4480
rect 10324 4437 10333 4471
rect 10333 4437 10367 4471
rect 10367 4437 10376 4471
rect 10324 4428 10376 4437
rect 22468 4428 22520 4480
rect 22836 4428 22888 4480
rect 3662 4326 3714 4378
rect 3726 4326 3778 4378
rect 3790 4326 3842 4378
rect 3854 4326 3906 4378
rect 3918 4326 3970 4378
rect 2320 4224 2372 4276
rect 2872 4224 2924 4276
rect 4436 4224 4488 4276
rect 4804 4224 4856 4276
rect 10232 4267 10284 4276
rect 10232 4233 10241 4267
rect 10241 4233 10275 4267
rect 10275 4233 10284 4267
rect 10232 4224 10284 4233
rect 10692 4224 10744 4276
rect 22836 4267 22888 4276
rect 22836 4233 22845 4267
rect 22845 4233 22879 4267
rect 22879 4233 22888 4267
rect 22836 4224 22888 4233
rect 1676 4131 1728 4140
rect 1676 4097 1685 4131
rect 1685 4097 1719 4131
rect 1719 4097 1728 4131
rect 1676 4088 1728 4097
rect 3240 4131 3292 4140
rect 3240 4097 3249 4131
rect 3249 4097 3283 4131
rect 3283 4097 3292 4131
rect 3240 4088 3292 4097
rect 4068 4156 4120 4208
rect 5632 4131 5684 4140
rect 5632 4097 5641 4131
rect 5641 4097 5675 4131
rect 5675 4097 5684 4131
rect 5632 4088 5684 4097
rect 11980 4088 12032 4140
rect 1768 4020 1820 4072
rect 3148 4020 3200 4072
rect 2964 3952 3016 4004
rect 4068 4063 4120 4072
rect 4068 4029 4077 4063
rect 4077 4029 4111 4063
rect 4111 4029 4120 4063
rect 4068 4020 4120 4029
rect 4344 4063 4396 4072
rect 4344 4029 4378 4063
rect 4378 4029 4396 4063
rect 4344 4020 4396 4029
rect 4804 4020 4856 4072
rect 4160 3952 4212 4004
rect 10232 4020 10284 4072
rect 11152 4063 11204 4072
rect 11152 4029 11161 4063
rect 11161 4029 11195 4063
rect 11195 4029 11204 4063
rect 11152 4020 11204 4029
rect 23020 4063 23072 4072
rect 23020 4029 23029 4063
rect 23029 4029 23063 4063
rect 23063 4029 23072 4063
rect 23020 4020 23072 4029
rect 10048 3952 10100 4004
rect 5448 3927 5500 3936
rect 5448 3893 5457 3927
rect 5457 3893 5491 3927
rect 5491 3893 5500 3927
rect 5448 3884 5500 3893
rect 9404 3884 9456 3936
rect 4322 3782 4374 3834
rect 4386 3782 4438 3834
rect 4450 3782 4502 3834
rect 4514 3782 4566 3834
rect 4578 3782 4630 3834
rect 3332 3680 3384 3732
rect 2964 3655 3016 3664
rect 2964 3621 2973 3655
rect 2973 3621 3007 3655
rect 3007 3621 3016 3655
rect 2964 3612 3016 3621
rect 3148 3655 3200 3664
rect 3148 3621 3157 3655
rect 3157 3621 3191 3655
rect 3191 3621 3200 3655
rect 4712 3723 4764 3732
rect 4712 3689 4721 3723
rect 4721 3689 4755 3723
rect 4755 3689 4764 3723
rect 4712 3680 4764 3689
rect 3148 3612 3200 3621
rect 3516 3655 3568 3664
rect 3516 3621 3550 3655
rect 3550 3621 3568 3655
rect 3516 3612 3568 3621
rect 4160 3612 4212 3664
rect 5448 3612 5500 3664
rect 2872 3587 2924 3596
rect 2872 3553 2881 3587
rect 2881 3553 2915 3587
rect 2915 3553 2924 3587
rect 2872 3544 2924 3553
rect 3056 3544 3108 3596
rect 4068 3544 4120 3596
rect 4804 3544 4856 3596
rect 3662 3238 3714 3290
rect 3726 3238 3778 3290
rect 3790 3238 3842 3290
rect 3854 3238 3906 3290
rect 3918 3238 3970 3290
rect 3424 3179 3476 3188
rect 3424 3145 3433 3179
rect 3433 3145 3467 3179
rect 3467 3145 3476 3179
rect 3424 3136 3476 3145
rect 2872 3000 2924 3052
rect 3148 2932 3200 2984
rect 4160 2932 4212 2984
rect 4322 2694 4374 2746
rect 4386 2694 4438 2746
rect 4450 2694 4502 2746
rect 4514 2694 4566 2746
rect 4578 2694 4630 2746
rect 3662 2150 3714 2202
rect 3726 2150 3778 2202
rect 3790 2150 3842 2202
rect 3854 2150 3906 2202
rect 3918 2150 3970 2202
rect 4322 1606 4374 1658
rect 4386 1606 4438 1658
rect 4450 1606 4502 1658
rect 4514 1606 4566 1658
rect 4578 1606 4630 1658
rect 3662 1062 3714 1114
rect 3726 1062 3778 1114
rect 3790 1062 3842 1114
rect 3854 1062 3906 1114
rect 3918 1062 3970 1114
rect 4322 518 4374 570
rect 4386 518 4438 570
rect 4450 518 4502 570
rect 4514 518 4566 570
rect 4578 518 4630 570
<< metal2 >>
rect 1674 23746 1730 24000
rect 4618 23746 4674 24000
rect 1674 23718 1808 23746
rect 1674 23600 1730 23718
rect 1780 23186 1808 23718
rect 4618 23718 4936 23746
rect 4618 23600 4674 23718
rect 4322 23420 4630 23429
rect 4322 23418 4328 23420
rect 4384 23418 4408 23420
rect 4464 23418 4488 23420
rect 4544 23418 4568 23420
rect 4624 23418 4630 23420
rect 4384 23366 4386 23418
rect 4566 23366 4568 23418
rect 4322 23364 4328 23366
rect 4384 23364 4408 23366
rect 4464 23364 4488 23366
rect 4544 23364 4568 23366
rect 4624 23364 4630 23366
rect 4322 23355 4630 23364
rect 4908 23254 4936 23718
rect 7562 23600 7618 24000
rect 10506 23600 10562 24000
rect 13450 23746 13506 24000
rect 16394 23746 16450 24000
rect 19338 23746 19394 24000
rect 13450 23718 13584 23746
rect 13450 23600 13506 23718
rect 5264 23316 5316 23322
rect 5264 23258 5316 23264
rect 3424 23248 3476 23254
rect 3424 23190 3476 23196
rect 4896 23248 4948 23254
rect 4896 23190 4948 23196
rect 1768 23180 1820 23186
rect 1768 23122 1820 23128
rect 2780 23180 2832 23186
rect 2780 23122 2832 23128
rect 2792 19922 2820 23122
rect 3436 23118 3464 23190
rect 5276 23186 5304 23258
rect 7576 23186 7604 23600
rect 10520 23254 10548 23600
rect 10508 23248 10560 23254
rect 10508 23190 10560 23196
rect 13556 23186 13584 23718
rect 16394 23718 16528 23746
rect 16394 23600 16450 23718
rect 16500 23186 16528 23718
rect 19338 23718 19472 23746
rect 19338 23600 19394 23718
rect 19444 23186 19472 23718
rect 22282 23600 22338 24000
rect 22296 23186 22324 23600
rect 4344 23180 4396 23186
rect 4344 23122 4396 23128
rect 4988 23180 5040 23186
rect 4988 23122 5040 23128
rect 5264 23180 5316 23186
rect 5264 23122 5316 23128
rect 7564 23180 7616 23186
rect 7564 23122 7616 23128
rect 13544 23180 13596 23186
rect 13544 23122 13596 23128
rect 16488 23180 16540 23186
rect 16488 23122 16540 23128
rect 17960 23180 18012 23186
rect 17960 23122 18012 23128
rect 18788 23180 18840 23186
rect 18788 23122 18840 23128
rect 19432 23180 19484 23186
rect 19432 23122 19484 23128
rect 22284 23180 22336 23186
rect 22284 23122 22336 23128
rect 3424 23112 3476 23118
rect 3424 23054 3476 23060
rect 2872 23044 2924 23050
rect 2872 22986 2924 22992
rect 2884 22438 2912 22986
rect 3056 22976 3108 22982
rect 3056 22918 3108 22924
rect 3068 22574 3096 22918
rect 3436 22574 3464 23054
rect 3662 22876 3970 22885
rect 3662 22874 3668 22876
rect 3724 22874 3748 22876
rect 3804 22874 3828 22876
rect 3884 22874 3908 22876
rect 3964 22874 3970 22876
rect 3724 22822 3726 22874
rect 3906 22822 3908 22874
rect 3662 22820 3668 22822
rect 3724 22820 3748 22822
rect 3804 22820 3828 22822
rect 3884 22820 3908 22822
rect 3964 22820 3970 22822
rect 3662 22811 3970 22820
rect 4356 22574 4384 23122
rect 4712 22772 4764 22778
rect 4712 22714 4764 22720
rect 4724 22574 4752 22714
rect 3056 22568 3108 22574
rect 3056 22510 3108 22516
rect 3424 22568 3476 22574
rect 3424 22510 3476 22516
rect 4344 22568 4396 22574
rect 4344 22510 4396 22516
rect 4712 22568 4764 22574
rect 4712 22510 4764 22516
rect 4804 22568 4856 22574
rect 4804 22510 4856 22516
rect 2872 22432 2924 22438
rect 2872 22374 2924 22380
rect 2884 19990 2912 22374
rect 2872 19984 2924 19990
rect 2872 19926 2924 19932
rect 3332 19984 3384 19990
rect 3332 19926 3384 19932
rect 2780 19916 2832 19922
rect 2780 19858 2832 19864
rect 2792 19310 2820 19858
rect 2884 19446 2912 19926
rect 3148 19712 3200 19718
rect 3148 19654 3200 19660
rect 3240 19712 3292 19718
rect 3240 19654 3292 19660
rect 3160 19446 3188 19654
rect 2872 19440 2924 19446
rect 2872 19382 2924 19388
rect 3148 19440 3200 19446
rect 3148 19382 3200 19388
rect 2780 19304 2832 19310
rect 2780 19246 2832 19252
rect 2792 18902 2820 19246
rect 2780 18896 2832 18902
rect 2780 18838 2832 18844
rect 2792 17814 2820 18838
rect 2780 17808 2832 17814
rect 2780 17750 2832 17756
rect 2884 16658 2912 19382
rect 3252 18698 3280 19654
rect 3344 19310 3372 19926
rect 3436 19922 3464 22510
rect 4322 22332 4630 22341
rect 4322 22330 4328 22332
rect 4384 22330 4408 22332
rect 4464 22330 4488 22332
rect 4544 22330 4568 22332
rect 4624 22330 4630 22332
rect 4384 22278 4386 22330
rect 4566 22278 4568 22330
rect 4322 22276 4328 22278
rect 4384 22276 4408 22278
rect 4464 22276 4488 22278
rect 4544 22276 4568 22278
rect 4624 22276 4630 22278
rect 4322 22267 4630 22276
rect 4252 22092 4304 22098
rect 4252 22034 4304 22040
rect 3662 21788 3970 21797
rect 3662 21786 3668 21788
rect 3724 21786 3748 21788
rect 3804 21786 3828 21788
rect 3884 21786 3908 21788
rect 3964 21786 3970 21788
rect 3724 21734 3726 21786
rect 3906 21734 3908 21786
rect 3662 21732 3668 21734
rect 3724 21732 3748 21734
rect 3804 21732 3828 21734
rect 3884 21732 3908 21734
rect 3964 21732 3970 21734
rect 3662 21723 3970 21732
rect 4264 21486 4292 22034
rect 4252 21480 4304 21486
rect 4252 21422 4304 21428
rect 3976 21344 4028 21350
rect 3976 21286 4028 21292
rect 3988 20890 4016 21286
rect 4264 21010 4292 21422
rect 4322 21244 4630 21253
rect 4322 21242 4328 21244
rect 4384 21242 4408 21244
rect 4464 21242 4488 21244
rect 4544 21242 4568 21244
rect 4624 21242 4630 21244
rect 4384 21190 4386 21242
rect 4566 21190 4568 21242
rect 4322 21188 4328 21190
rect 4384 21188 4408 21190
rect 4464 21188 4488 21190
rect 4544 21188 4568 21190
rect 4624 21188 4630 21190
rect 4322 21179 4630 21188
rect 4528 21072 4580 21078
rect 4724 21026 4752 22510
rect 4816 21486 4844 22510
rect 4804 21480 4856 21486
rect 4804 21422 4856 21428
rect 4528 21014 4580 21020
rect 4252 21004 4304 21010
rect 4252 20946 4304 20952
rect 3988 20862 4108 20890
rect 3662 20700 3970 20709
rect 3662 20698 3668 20700
rect 3724 20698 3748 20700
rect 3804 20698 3828 20700
rect 3884 20698 3908 20700
rect 3964 20698 3970 20700
rect 3724 20646 3726 20698
rect 3906 20646 3908 20698
rect 3662 20644 3668 20646
rect 3724 20644 3748 20646
rect 3804 20644 3828 20646
rect 3884 20644 3908 20646
rect 3964 20644 3970 20646
rect 3662 20635 3970 20644
rect 4080 20330 4108 20862
rect 4540 20602 4568 21014
rect 4632 20998 4752 21026
rect 4528 20596 4580 20602
rect 4528 20538 4580 20544
rect 4632 20398 4660 20998
rect 4804 20528 4856 20534
rect 4804 20470 4856 20476
rect 4620 20392 4672 20398
rect 4620 20334 4672 20340
rect 4068 20324 4120 20330
rect 4068 20266 4120 20272
rect 4080 19990 4108 20266
rect 4322 20156 4630 20165
rect 4322 20154 4328 20156
rect 4384 20154 4408 20156
rect 4464 20154 4488 20156
rect 4544 20154 4568 20156
rect 4624 20154 4630 20156
rect 4384 20102 4386 20154
rect 4566 20102 4568 20154
rect 4322 20100 4328 20102
rect 4384 20100 4408 20102
rect 4464 20100 4488 20102
rect 4544 20100 4568 20102
rect 4624 20100 4630 20102
rect 4322 20091 4630 20100
rect 4068 19984 4120 19990
rect 4068 19926 4120 19932
rect 3424 19916 3476 19922
rect 3424 19858 3476 19864
rect 3662 19612 3970 19621
rect 3662 19610 3668 19612
rect 3724 19610 3748 19612
rect 3804 19610 3828 19612
rect 3884 19610 3908 19612
rect 3964 19610 3970 19612
rect 3724 19558 3726 19610
rect 3906 19558 3908 19610
rect 3662 19556 3668 19558
rect 3724 19556 3748 19558
rect 3804 19556 3828 19558
rect 3884 19556 3908 19558
rect 3964 19556 3970 19558
rect 3662 19547 3970 19556
rect 3700 19440 3752 19446
rect 3700 19382 3752 19388
rect 3332 19304 3384 19310
rect 3332 19246 3384 19252
rect 3608 19304 3660 19310
rect 3608 19246 3660 19252
rect 3240 18692 3292 18698
rect 3240 18634 3292 18640
rect 3252 17728 3280 18634
rect 3344 18290 3372 19246
rect 3516 19236 3568 19242
rect 3516 19178 3568 19184
rect 3528 18630 3556 19178
rect 3620 18970 3648 19246
rect 3608 18964 3660 18970
rect 3608 18906 3660 18912
rect 3712 18834 3740 19382
rect 4252 19168 4304 19174
rect 4252 19110 4304 19116
rect 3700 18828 3752 18834
rect 3700 18770 3752 18776
rect 4160 18828 4212 18834
rect 4160 18770 4212 18776
rect 3516 18624 3568 18630
rect 3516 18566 3568 18572
rect 4068 18624 4120 18630
rect 4068 18566 4120 18572
rect 3662 18524 3970 18533
rect 3662 18522 3668 18524
rect 3724 18522 3748 18524
rect 3804 18522 3828 18524
rect 3884 18522 3908 18524
rect 3964 18522 3970 18524
rect 3724 18470 3726 18522
rect 3906 18470 3908 18522
rect 3662 18468 3668 18470
rect 3724 18468 3748 18470
rect 3804 18468 3828 18470
rect 3884 18468 3908 18470
rect 3964 18468 3970 18470
rect 3662 18459 3970 18468
rect 3332 18284 3384 18290
rect 3332 18226 3384 18232
rect 3424 17808 3476 17814
rect 3424 17750 3476 17756
rect 3332 17740 3384 17746
rect 3252 17700 3332 17728
rect 3332 17682 3384 17688
rect 3148 17672 3200 17678
rect 3148 17614 3200 17620
rect 3160 16658 3188 17614
rect 3344 17066 3372 17682
rect 3332 17060 3384 17066
rect 3332 17002 3384 17008
rect 3436 16998 3464 17750
rect 3662 17436 3970 17445
rect 3662 17434 3668 17436
rect 3724 17434 3748 17436
rect 3804 17434 3828 17436
rect 3884 17434 3908 17436
rect 3964 17434 3970 17436
rect 3724 17382 3726 17434
rect 3906 17382 3908 17434
rect 3662 17380 3668 17382
rect 3724 17380 3748 17382
rect 3804 17380 3828 17382
rect 3884 17380 3908 17382
rect 3964 17380 3970 17382
rect 3662 17371 3970 17380
rect 3516 17332 3568 17338
rect 3516 17274 3568 17280
rect 3424 16992 3476 16998
rect 3424 16934 3476 16940
rect 2872 16652 2924 16658
rect 2872 16594 2924 16600
rect 3148 16652 3200 16658
rect 3148 16594 3200 16600
rect 2884 16130 2912 16594
rect 3056 16584 3108 16590
rect 3056 16526 3108 16532
rect 2792 16102 3004 16130
rect 2792 14482 2820 16102
rect 2976 15978 3004 16102
rect 2872 15972 2924 15978
rect 2872 15914 2924 15920
rect 2964 15972 3016 15978
rect 2964 15914 3016 15920
rect 2884 14482 2912 15914
rect 3068 15910 3096 16526
rect 3160 16182 3188 16594
rect 3148 16176 3200 16182
rect 3148 16118 3200 16124
rect 3056 15904 3108 15910
rect 3056 15846 3108 15852
rect 3068 15706 3096 15846
rect 3056 15700 3108 15706
rect 3056 15642 3108 15648
rect 3160 15570 3188 16118
rect 3436 16114 3464 16934
rect 3528 16658 3556 17274
rect 4080 17218 4108 18566
rect 3896 17190 4108 17218
rect 3608 17060 3660 17066
rect 3608 17002 3660 17008
rect 3516 16652 3568 16658
rect 3516 16594 3568 16600
rect 3620 16538 3648 17002
rect 3896 16658 3924 17190
rect 4068 16992 4120 16998
rect 4068 16934 4120 16940
rect 4080 16658 4108 16934
rect 4172 16794 4200 18770
rect 4264 18408 4292 19110
rect 4322 19068 4630 19077
rect 4322 19066 4328 19068
rect 4384 19066 4408 19068
rect 4464 19066 4488 19068
rect 4544 19066 4568 19068
rect 4624 19066 4630 19068
rect 4384 19014 4386 19066
rect 4566 19014 4568 19066
rect 4322 19012 4328 19014
rect 4384 19012 4408 19014
rect 4464 19012 4488 19014
rect 4544 19012 4568 19014
rect 4624 19012 4630 19014
rect 4322 19003 4630 19012
rect 4264 18380 4384 18408
rect 4252 18284 4304 18290
rect 4252 18226 4304 18232
rect 4160 16788 4212 16794
rect 4160 16730 4212 16736
rect 3884 16652 3936 16658
rect 3884 16594 3936 16600
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 3528 16522 3648 16538
rect 3516 16516 3648 16522
rect 3568 16510 3648 16516
rect 3516 16458 3568 16464
rect 3424 16108 3476 16114
rect 3424 16050 3476 16056
rect 3528 16046 3556 16458
rect 3662 16348 3970 16357
rect 3662 16346 3668 16348
rect 3724 16346 3748 16348
rect 3804 16346 3828 16348
rect 3884 16346 3908 16348
rect 3964 16346 3970 16348
rect 3724 16294 3726 16346
rect 3906 16294 3908 16346
rect 3662 16292 3668 16294
rect 3724 16292 3748 16294
rect 3804 16292 3828 16294
rect 3884 16292 3908 16294
rect 3964 16292 3970 16294
rect 3662 16283 3970 16292
rect 4172 16114 4200 16730
rect 3976 16108 4028 16114
rect 3976 16050 4028 16056
rect 4160 16108 4212 16114
rect 4160 16050 4212 16056
rect 3516 16040 3568 16046
rect 3516 15982 3568 15988
rect 3608 15972 3660 15978
rect 3608 15914 3660 15920
rect 3700 15972 3752 15978
rect 3700 15914 3752 15920
rect 3148 15564 3200 15570
rect 3148 15506 3200 15512
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 3620 15450 3648 15914
rect 3712 15638 3740 15914
rect 3792 15904 3844 15910
rect 3792 15846 3844 15852
rect 3804 15638 3832 15846
rect 3700 15632 3752 15638
rect 3700 15574 3752 15580
rect 3792 15632 3844 15638
rect 3792 15574 3844 15580
rect 3988 15570 4016 16050
rect 4264 15858 4292 18226
rect 4356 18222 4384 18380
rect 4344 18216 4396 18222
rect 4344 18158 4396 18164
rect 4322 17980 4630 17989
rect 4322 17978 4328 17980
rect 4384 17978 4408 17980
rect 4464 17978 4488 17980
rect 4544 17978 4568 17980
rect 4624 17978 4630 17980
rect 4384 17926 4386 17978
rect 4566 17926 4568 17978
rect 4322 17924 4328 17926
rect 4384 17924 4408 17926
rect 4464 17924 4488 17926
rect 4544 17924 4568 17926
rect 4624 17924 4630 17926
rect 4322 17915 4630 17924
rect 4322 16892 4630 16901
rect 4322 16890 4328 16892
rect 4384 16890 4408 16892
rect 4464 16890 4488 16892
rect 4544 16890 4568 16892
rect 4624 16890 4630 16892
rect 4384 16838 4386 16890
rect 4566 16838 4568 16890
rect 4322 16836 4328 16838
rect 4384 16836 4408 16838
rect 4464 16836 4488 16838
rect 4544 16836 4568 16838
rect 4624 16836 4630 16838
rect 4322 16827 4630 16836
rect 4620 16584 4672 16590
rect 4620 16526 4672 16532
rect 4632 16046 4660 16526
rect 4620 16040 4672 16046
rect 4672 16000 4752 16028
rect 4620 15982 4672 15988
rect 4172 15830 4292 15858
rect 3884 15564 3936 15570
rect 3884 15506 3936 15512
rect 3976 15564 4028 15570
rect 3976 15506 4028 15512
rect 3896 15450 3924 15506
rect 2976 14618 3004 15438
rect 3620 15422 3924 15450
rect 3662 15260 3970 15269
rect 3662 15258 3668 15260
rect 3724 15258 3748 15260
rect 3804 15258 3828 15260
rect 3884 15258 3908 15260
rect 3964 15258 3970 15260
rect 3724 15206 3726 15258
rect 3906 15206 3908 15258
rect 3662 15204 3668 15206
rect 3724 15204 3748 15206
rect 3804 15204 3828 15206
rect 3884 15204 3908 15206
rect 3964 15204 3970 15206
rect 3662 15195 3970 15204
rect 4172 14958 4200 15830
rect 4322 15804 4630 15813
rect 4322 15802 4328 15804
rect 4384 15802 4408 15804
rect 4464 15802 4488 15804
rect 4544 15802 4568 15804
rect 4624 15802 4630 15804
rect 4384 15750 4386 15802
rect 4566 15750 4568 15802
rect 4322 15748 4328 15750
rect 4384 15748 4408 15750
rect 4464 15748 4488 15750
rect 4544 15748 4568 15750
rect 4624 15748 4630 15750
rect 4322 15739 4630 15748
rect 4724 15570 4752 16000
rect 4712 15564 4764 15570
rect 4712 15506 4764 15512
rect 4712 15428 4764 15434
rect 4712 15370 4764 15376
rect 4252 15360 4304 15366
rect 4252 15302 4304 15308
rect 4264 15026 4292 15302
rect 4724 15026 4752 15370
rect 4252 15020 4304 15026
rect 4252 14962 4304 14968
rect 4712 15020 4764 15026
rect 4712 14962 4764 14968
rect 4160 14952 4212 14958
rect 4160 14894 4212 14900
rect 2964 14612 3016 14618
rect 2964 14554 3016 14560
rect 3424 14612 3476 14618
rect 3424 14554 3476 14560
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 2872 14476 2924 14482
rect 2872 14418 2924 14424
rect 2792 13870 2820 14418
rect 2884 13870 2912 14418
rect 3148 13932 3200 13938
rect 3148 13874 3200 13880
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2872 13864 2924 13870
rect 2872 13806 2924 13812
rect 2792 12442 2820 13806
rect 3160 13802 3188 13874
rect 3436 13870 3464 14554
rect 4172 14550 4200 14894
rect 4160 14544 4212 14550
rect 4160 14486 4212 14492
rect 4264 14482 4292 14962
rect 4322 14716 4630 14725
rect 4322 14714 4328 14716
rect 4384 14714 4408 14716
rect 4464 14714 4488 14716
rect 4544 14714 4568 14716
rect 4624 14714 4630 14716
rect 4384 14662 4386 14714
rect 4566 14662 4568 14714
rect 4322 14660 4328 14662
rect 4384 14660 4408 14662
rect 4464 14660 4488 14662
rect 4544 14660 4568 14662
rect 4624 14660 4630 14662
rect 4322 14651 4630 14660
rect 4252 14476 4304 14482
rect 4252 14418 4304 14424
rect 3662 14172 3970 14181
rect 3662 14170 3668 14172
rect 3724 14170 3748 14172
rect 3804 14170 3828 14172
rect 3884 14170 3908 14172
rect 3964 14170 3970 14172
rect 3724 14118 3726 14170
rect 3906 14118 3908 14170
rect 3662 14116 3668 14118
rect 3724 14116 3748 14118
rect 3804 14116 3828 14118
rect 3884 14116 3908 14118
rect 3964 14116 3970 14118
rect 3662 14107 3970 14116
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 3148 13796 3200 13802
rect 3148 13738 3200 13744
rect 3516 13796 3568 13802
rect 3516 13738 3568 13744
rect 2780 12436 2832 12442
rect 3160 12434 3188 13738
rect 3528 13274 3556 13738
rect 3792 13728 3844 13734
rect 3792 13670 3844 13676
rect 3804 13462 3832 13670
rect 4322 13628 4630 13637
rect 4322 13626 4328 13628
rect 4384 13626 4408 13628
rect 4464 13626 4488 13628
rect 4544 13626 4568 13628
rect 4624 13626 4630 13628
rect 4384 13574 4386 13626
rect 4566 13574 4568 13626
rect 4322 13572 4328 13574
rect 4384 13572 4408 13574
rect 4464 13572 4488 13574
rect 4544 13572 4568 13574
rect 4624 13572 4630 13574
rect 4322 13563 4630 13572
rect 3792 13456 3844 13462
rect 3792 13398 3844 13404
rect 3436 13246 3556 13274
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 3436 13190 3464 13246
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 3436 12434 3464 13126
rect 3662 13084 3970 13093
rect 3662 13082 3668 13084
rect 3724 13082 3748 13084
rect 3804 13082 3828 13084
rect 3884 13082 3908 13084
rect 3964 13082 3970 13084
rect 3724 13030 3726 13082
rect 3906 13030 3908 13082
rect 3662 13028 3668 13030
rect 3724 13028 3748 13030
rect 3804 13028 3828 13030
rect 3884 13028 3908 13030
rect 3964 13028 3970 13030
rect 3662 13019 3970 13028
rect 4252 12640 4304 12646
rect 4252 12582 4304 12588
rect 3160 12406 3280 12434
rect 3436 12406 3556 12434
rect 2780 12378 2832 12384
rect 3252 12238 3280 12406
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3332 12232 3384 12238
rect 3332 12174 3384 12180
rect 3252 11626 3280 12174
rect 3344 11898 3372 12174
rect 3332 11892 3384 11898
rect 3332 11834 3384 11840
rect 3240 11620 3292 11626
rect 3240 11562 3292 11568
rect 3240 11144 3292 11150
rect 3240 11086 3292 11092
rect 3056 9036 3108 9042
rect 3056 8978 3108 8984
rect 3068 8022 3096 8978
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 3160 8430 3188 8774
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 3148 8084 3200 8090
rect 3148 8026 3200 8032
rect 3056 8016 3108 8022
rect 3056 7958 3108 7964
rect 3160 7954 3188 8026
rect 3148 7948 3200 7954
rect 3148 7890 3200 7896
rect 2320 7744 2372 7750
rect 2320 7686 2372 7692
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2136 7268 2188 7274
rect 2136 7210 2188 7216
rect 2148 7002 2176 7210
rect 2136 6996 2188 7002
rect 2136 6938 2188 6944
rect 2332 6662 2360 7686
rect 2424 7002 2452 7686
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 2412 6996 2464 7002
rect 2412 6938 2464 6944
rect 2780 6928 2832 6934
rect 2780 6870 2832 6876
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 2792 5370 2820 6870
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 2504 5024 2556 5030
rect 2504 4966 2556 4972
rect 2516 4758 2544 4966
rect 2504 4752 2556 4758
rect 2504 4694 2556 4700
rect 1676 4684 1728 4690
rect 1676 4626 1728 4632
rect 1688 4146 1716 4626
rect 2320 4616 2372 4622
rect 2320 4558 2372 4564
rect 1768 4480 1820 4486
rect 1768 4422 1820 4428
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 1780 4078 1808 4422
rect 2332 4282 2360 4558
rect 2792 4486 2820 5306
rect 2884 5166 2912 7346
rect 2976 6662 3004 7686
rect 3160 7546 3188 7890
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 3160 7290 3188 7482
rect 3252 7410 3280 11086
rect 3344 10130 3372 11834
rect 3332 10124 3384 10130
rect 3332 10066 3384 10072
rect 3344 9042 3372 10066
rect 3528 10062 3556 12406
rect 4264 12374 4292 12582
rect 4322 12540 4630 12549
rect 4322 12538 4328 12540
rect 4384 12538 4408 12540
rect 4464 12538 4488 12540
rect 4544 12538 4568 12540
rect 4624 12538 4630 12540
rect 4384 12486 4386 12538
rect 4566 12486 4568 12538
rect 4322 12484 4328 12486
rect 4384 12484 4408 12486
rect 4464 12484 4488 12486
rect 4544 12484 4568 12486
rect 4624 12484 4630 12486
rect 4322 12475 4630 12484
rect 4252 12368 4304 12374
rect 4252 12310 4304 12316
rect 4620 12300 4672 12306
rect 4724 12288 4752 13262
rect 4816 12646 4844 20470
rect 5000 20398 5028 23122
rect 5816 23112 5868 23118
rect 5816 23054 5868 23060
rect 13912 23112 13964 23118
rect 13912 23054 13964 23060
rect 15200 23112 15252 23118
rect 15200 23054 15252 23060
rect 15476 23112 15528 23118
rect 15476 23054 15528 23060
rect 5080 22500 5132 22506
rect 5080 22442 5132 22448
rect 5092 22098 5120 22442
rect 5828 22098 5856 23054
rect 7288 23044 7340 23050
rect 7288 22986 7340 22992
rect 7196 22976 7248 22982
rect 7196 22918 7248 22924
rect 7208 22778 7236 22918
rect 7300 22778 7328 22986
rect 9588 22976 9640 22982
rect 9588 22918 9640 22924
rect 7196 22772 7248 22778
rect 7196 22714 7248 22720
rect 7288 22772 7340 22778
rect 7288 22714 7340 22720
rect 8208 22772 8260 22778
rect 8208 22714 8260 22720
rect 6000 22704 6052 22710
rect 6000 22646 6052 22652
rect 6012 22098 6040 22646
rect 6276 22568 6328 22574
rect 6276 22510 6328 22516
rect 6288 22166 6316 22510
rect 7104 22432 7156 22438
rect 7104 22374 7156 22380
rect 6828 22228 6880 22234
rect 6828 22170 6880 22176
rect 6276 22160 6328 22166
rect 6276 22102 6328 22108
rect 6840 22114 6868 22170
rect 5080 22092 5132 22098
rect 5080 22034 5132 22040
rect 5816 22092 5868 22098
rect 5816 22034 5868 22040
rect 6000 22092 6052 22098
rect 6000 22034 6052 22040
rect 5092 21010 5120 22034
rect 5172 21956 5224 21962
rect 5172 21898 5224 21904
rect 5184 21554 5212 21898
rect 5908 21888 5960 21894
rect 5908 21830 5960 21836
rect 5172 21548 5224 21554
rect 5172 21490 5224 21496
rect 5080 21004 5132 21010
rect 5080 20946 5132 20952
rect 4988 20392 5040 20398
rect 4988 20334 5040 20340
rect 4896 20324 4948 20330
rect 4896 20266 4948 20272
rect 4908 19922 4936 20266
rect 5000 20074 5028 20334
rect 5000 20058 5120 20074
rect 5000 20052 5132 20058
rect 5000 20046 5080 20052
rect 5080 19994 5132 20000
rect 4988 19984 5040 19990
rect 4988 19926 5040 19932
rect 4896 19916 4948 19922
rect 4896 19858 4948 19864
rect 4896 19780 4948 19786
rect 4896 19722 4948 19728
rect 4908 19378 4936 19722
rect 4896 19372 4948 19378
rect 4896 19314 4948 19320
rect 4908 18698 4936 19314
rect 5000 19310 5028 19926
rect 4988 19304 5040 19310
rect 4988 19246 5040 19252
rect 5184 19122 5212 21490
rect 5920 21486 5948 21830
rect 6288 21554 6316 22102
rect 6840 22094 6960 22114
rect 7116 22098 7144 22374
rect 7012 22094 7064 22098
rect 6840 22092 7064 22094
rect 6840 22086 7012 22092
rect 6368 21888 6420 21894
rect 6368 21830 6420 21836
rect 6276 21548 6328 21554
rect 6276 21490 6328 21496
rect 5908 21480 5960 21486
rect 5908 21422 5960 21428
rect 5908 21344 5960 21350
rect 5906 21312 5908 21321
rect 6184 21344 6236 21350
rect 5960 21312 5962 21321
rect 6184 21286 6236 21292
rect 5906 21247 5962 21256
rect 5264 20596 5316 20602
rect 5264 20538 5316 20544
rect 5276 20398 5304 20538
rect 5264 20392 5316 20398
rect 5264 20334 5316 20340
rect 5540 20392 5592 20398
rect 5540 20334 5592 20340
rect 5000 19094 5212 19122
rect 5000 18834 5028 19094
rect 5276 18970 5304 20334
rect 5448 19508 5500 19514
rect 5448 19450 5500 19456
rect 5264 18964 5316 18970
rect 5264 18906 5316 18912
rect 4988 18828 5040 18834
rect 4988 18770 5040 18776
rect 4896 18692 4948 18698
rect 4896 18634 4948 18640
rect 4896 18216 4948 18222
rect 4896 18158 4948 18164
rect 4804 12640 4856 12646
rect 4804 12582 4856 12588
rect 4672 12260 4752 12288
rect 4620 12242 4672 12248
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 3662 11996 3970 12005
rect 3662 11994 3668 11996
rect 3724 11994 3748 11996
rect 3804 11994 3828 11996
rect 3884 11994 3908 11996
rect 3964 11994 3970 11996
rect 3724 11942 3726 11994
rect 3906 11942 3908 11994
rect 3662 11940 3668 11942
rect 3724 11940 3748 11942
rect 3804 11940 3828 11942
rect 3884 11940 3908 11942
rect 3964 11940 3970 11942
rect 3662 11931 3970 11940
rect 4356 11694 4384 12038
rect 4632 11762 4660 12242
rect 4908 11762 4936 18158
rect 5000 14958 5028 18770
rect 5080 18760 5132 18766
rect 5080 18702 5132 18708
rect 5092 18154 5120 18702
rect 5276 18222 5304 18906
rect 5460 18766 5488 19450
rect 5552 18902 5580 20334
rect 6000 19712 6052 19718
rect 6000 19654 6052 19660
rect 6012 19310 6040 19654
rect 6000 19304 6052 19310
rect 6000 19246 6052 19252
rect 5540 18896 5592 18902
rect 5540 18838 5592 18844
rect 5448 18760 5500 18766
rect 5448 18702 5500 18708
rect 5264 18216 5316 18222
rect 5264 18158 5316 18164
rect 5080 18148 5132 18154
rect 5080 18090 5132 18096
rect 5092 17882 5120 18090
rect 5080 17876 5132 17882
rect 5080 17818 5132 17824
rect 5276 16658 5304 18158
rect 5448 17128 5500 17134
rect 5448 17070 5500 17076
rect 6092 17128 6144 17134
rect 6092 17070 6144 17076
rect 5460 16794 5488 17070
rect 5448 16788 5500 16794
rect 5448 16730 5500 16736
rect 5264 16652 5316 16658
rect 5264 16594 5316 16600
rect 5460 16046 5488 16730
rect 6104 16114 6132 17070
rect 6092 16108 6144 16114
rect 6092 16050 6144 16056
rect 5448 16040 5500 16046
rect 5448 15982 5500 15988
rect 4988 14952 5040 14958
rect 4988 14894 5040 14900
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5184 14482 5212 14758
rect 5368 14618 5396 14758
rect 5356 14612 5408 14618
rect 5356 14554 5408 14560
rect 5172 14476 5224 14482
rect 5172 14418 5224 14424
rect 5184 14006 5212 14418
rect 5460 14414 5488 15982
rect 5908 15020 5960 15026
rect 5908 14962 5960 14968
rect 5920 14414 5948 14962
rect 6092 14476 6144 14482
rect 6092 14418 6144 14424
rect 5448 14408 5500 14414
rect 5448 14350 5500 14356
rect 5908 14408 5960 14414
rect 5908 14350 5960 14356
rect 5172 14000 5224 14006
rect 5172 13942 5224 13948
rect 5460 13938 5488 14350
rect 6000 14340 6052 14346
rect 6000 14282 6052 14288
rect 6012 13938 6040 14282
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 6000 13932 6052 13938
rect 6000 13874 6052 13880
rect 5724 13728 5776 13734
rect 5724 13670 5776 13676
rect 5736 13462 5764 13670
rect 5724 13456 5776 13462
rect 5724 13398 5776 13404
rect 6012 13394 6040 13874
rect 6104 13870 6132 14418
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 6000 13388 6052 13394
rect 6000 13330 6052 13336
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 4988 12776 5040 12782
rect 4988 12718 5040 12724
rect 4620 11756 4672 11762
rect 4620 11698 4672 11704
rect 4896 11756 4948 11762
rect 4896 11698 4948 11704
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 4322 11452 4630 11461
rect 4322 11450 4328 11452
rect 4384 11450 4408 11452
rect 4464 11450 4488 11452
rect 4544 11450 4568 11452
rect 4624 11450 4630 11452
rect 4384 11398 4386 11450
rect 4566 11398 4568 11450
rect 4322 11396 4328 11398
rect 4384 11396 4408 11398
rect 4464 11396 4488 11398
rect 4544 11396 4568 11398
rect 4624 11396 4630 11398
rect 4322 11387 4630 11396
rect 4724 11286 4752 11494
rect 4712 11280 4764 11286
rect 4712 11222 4764 11228
rect 3662 10908 3970 10917
rect 3662 10906 3668 10908
rect 3724 10906 3748 10908
rect 3804 10906 3828 10908
rect 3884 10906 3908 10908
rect 3964 10906 3970 10908
rect 3724 10854 3726 10906
rect 3906 10854 3908 10906
rect 3662 10852 3668 10854
rect 3724 10852 3748 10854
rect 3804 10852 3828 10854
rect 3884 10852 3908 10854
rect 3964 10852 3970 10854
rect 3662 10843 3970 10852
rect 4322 10364 4630 10373
rect 4322 10362 4328 10364
rect 4384 10362 4408 10364
rect 4464 10362 4488 10364
rect 4544 10362 4568 10364
rect 4624 10362 4630 10364
rect 4384 10310 4386 10362
rect 4566 10310 4568 10362
rect 4322 10308 4328 10310
rect 4384 10308 4408 10310
rect 4464 10308 4488 10310
rect 4544 10308 4568 10310
rect 4624 10308 4630 10310
rect 4322 10299 4630 10308
rect 4896 10124 4948 10130
rect 4896 10066 4948 10072
rect 3516 10056 3568 10062
rect 3516 9998 3568 10004
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 4620 9920 4672 9926
rect 4620 9862 4672 9868
rect 3662 9820 3970 9829
rect 3662 9818 3668 9820
rect 3724 9818 3748 9820
rect 3804 9818 3828 9820
rect 3884 9818 3908 9820
rect 3964 9818 3970 9820
rect 3724 9766 3726 9818
rect 3906 9766 3908 9818
rect 3662 9764 3668 9766
rect 3724 9764 3748 9766
rect 3804 9764 3828 9766
rect 3884 9764 3908 9766
rect 3964 9764 3970 9766
rect 3662 9755 3970 9764
rect 3332 9036 3384 9042
rect 3332 8978 3384 8984
rect 4080 8974 4108 9862
rect 4632 9722 4660 9862
rect 4620 9716 4672 9722
rect 4620 9658 4672 9664
rect 4724 9586 4752 9998
rect 4804 9988 4856 9994
rect 4804 9930 4856 9936
rect 4816 9586 4844 9930
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 4804 9580 4856 9586
rect 4804 9522 4856 9528
rect 4712 9444 4764 9450
rect 4712 9386 4764 9392
rect 4322 9276 4630 9285
rect 4322 9274 4328 9276
rect 4384 9274 4408 9276
rect 4464 9274 4488 9276
rect 4544 9274 4568 9276
rect 4624 9274 4630 9276
rect 4384 9222 4386 9274
rect 4566 9222 4568 9274
rect 4322 9220 4328 9222
rect 4384 9220 4408 9222
rect 4464 9220 4488 9222
rect 4544 9220 4568 9222
rect 4624 9220 4630 9222
rect 4322 9211 4630 9220
rect 4160 9036 4212 9042
rect 4160 8978 4212 8984
rect 3516 8968 3568 8974
rect 3516 8910 3568 8916
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 3424 8356 3476 8362
rect 3424 8298 3476 8304
rect 3436 7954 3464 8298
rect 3528 8090 3556 8910
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 3662 8732 3970 8741
rect 3662 8730 3668 8732
rect 3724 8730 3748 8732
rect 3804 8730 3828 8732
rect 3884 8730 3908 8732
rect 3964 8730 3970 8732
rect 3724 8678 3726 8730
rect 3906 8678 3908 8730
rect 3662 8676 3668 8678
rect 3724 8676 3748 8678
rect 3804 8676 3828 8678
rect 3884 8676 3908 8678
rect 3964 8676 3970 8678
rect 3662 8667 3970 8676
rect 4080 8634 4108 8774
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 4172 8362 4200 8978
rect 4724 8362 4752 9386
rect 4816 8362 4844 9522
rect 4908 9518 4936 10066
rect 5000 9654 5028 12718
rect 5276 11762 5304 12786
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 5368 12442 5396 12718
rect 5356 12436 5408 12442
rect 5356 12378 5408 12384
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 5092 11354 5120 11494
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 5092 10062 5120 11290
rect 5276 11150 5304 11698
rect 6196 11354 6224 21286
rect 6288 20466 6316 21490
rect 6380 21350 6408 21830
rect 6840 21554 6868 22086
rect 6932 22066 7012 22086
rect 7012 22034 7064 22040
rect 7104 22092 7156 22098
rect 7300 22094 7328 22714
rect 7472 22568 7524 22574
rect 7472 22510 7524 22516
rect 7840 22568 7892 22574
rect 7840 22510 7892 22516
rect 7300 22066 7420 22094
rect 7104 22034 7156 22040
rect 6920 22024 6972 22030
rect 6920 21966 6972 21972
rect 6932 21690 6960 21966
rect 6920 21684 6972 21690
rect 6920 21626 6972 21632
rect 6828 21548 6880 21554
rect 6828 21490 6880 21496
rect 6368 21344 6420 21350
rect 6368 21286 6420 21292
rect 6380 20942 6408 21286
rect 7116 21078 7144 22034
rect 7194 21992 7250 22001
rect 7194 21927 7250 21936
rect 7104 21072 7156 21078
rect 7104 21014 7156 21020
rect 7208 21010 7236 21927
rect 7288 21888 7340 21894
rect 7286 21856 7288 21865
rect 7340 21856 7342 21865
rect 7286 21791 7342 21800
rect 7392 21010 7420 22066
rect 7484 21486 7512 22510
rect 7748 22500 7800 22506
rect 7748 22442 7800 22448
rect 7760 22098 7788 22442
rect 7748 22092 7800 22098
rect 7748 22034 7800 22040
rect 7760 21690 7788 22034
rect 7748 21684 7800 21690
rect 7748 21626 7800 21632
rect 7564 21616 7616 21622
rect 7564 21558 7616 21564
rect 7472 21480 7524 21486
rect 7472 21422 7524 21428
rect 7576 21010 7604 21558
rect 7852 21554 7880 22510
rect 8220 22438 8248 22714
rect 8484 22568 8536 22574
rect 8484 22510 8536 22516
rect 7932 22432 7984 22438
rect 7932 22374 7984 22380
rect 8208 22432 8260 22438
rect 8208 22374 8260 22380
rect 7944 22098 7972 22374
rect 8496 22234 8524 22510
rect 8668 22432 8720 22438
rect 8668 22374 8720 22380
rect 8484 22228 8536 22234
rect 8484 22170 8536 22176
rect 8116 22160 8168 22166
rect 8116 22102 8168 22108
rect 7932 22092 7984 22098
rect 7932 22034 7984 22040
rect 8128 21690 8156 22102
rect 8300 22092 8352 22098
rect 8496 22094 8524 22170
rect 8680 22098 8708 22374
rect 8300 22034 8352 22040
rect 8404 22066 8524 22094
rect 8576 22092 8628 22098
rect 8116 21684 8168 21690
rect 8116 21626 8168 21632
rect 8312 21622 8340 22034
rect 8300 21616 8352 21622
rect 8300 21558 8352 21564
rect 7840 21548 7892 21554
rect 7840 21490 7892 21496
rect 7656 21480 7708 21486
rect 7656 21422 7708 21428
rect 7668 21332 7696 21422
rect 8208 21412 8260 21418
rect 8208 21354 8260 21360
rect 7748 21344 7800 21350
rect 7668 21304 7748 21332
rect 7748 21286 7800 21292
rect 8220 21010 8248 21354
rect 7196 21004 7248 21010
rect 7196 20946 7248 20952
rect 7380 21004 7432 21010
rect 7380 20946 7432 20952
rect 7564 21004 7616 21010
rect 7564 20946 7616 20952
rect 8208 21004 8260 21010
rect 8208 20946 8260 20952
rect 6368 20936 6420 20942
rect 6368 20878 6420 20884
rect 7208 20754 7236 20946
rect 7116 20726 7236 20754
rect 6276 20460 6328 20466
rect 6276 20402 6328 20408
rect 6736 20256 6788 20262
rect 6736 20198 6788 20204
rect 6748 19378 6776 20198
rect 6736 19372 6788 19378
rect 6736 19314 6788 19320
rect 6276 19168 6328 19174
rect 6276 19110 6328 19116
rect 6288 18902 6316 19110
rect 6276 18896 6328 18902
rect 6276 18838 6328 18844
rect 6288 18426 6316 18838
rect 6644 18828 6696 18834
rect 6748 18816 6776 19314
rect 7116 19174 7144 20726
rect 7392 20398 7420 20946
rect 7380 20392 7432 20398
rect 7380 20334 7432 20340
rect 7392 19938 7420 20334
rect 7392 19910 7512 19938
rect 7196 19440 7248 19446
rect 7196 19382 7248 19388
rect 7104 19168 7156 19174
rect 7104 19110 7156 19116
rect 6696 18788 6776 18816
rect 6840 18788 7052 18816
rect 6644 18770 6696 18776
rect 6840 18698 6868 18788
rect 6828 18692 6880 18698
rect 6828 18634 6880 18640
rect 6920 18692 6972 18698
rect 6920 18634 6972 18640
rect 6276 18420 6328 18426
rect 6276 18362 6328 18368
rect 6276 16652 6328 16658
rect 6276 16594 6328 16600
rect 6288 16046 6316 16594
rect 6460 16584 6512 16590
rect 6460 16526 6512 16532
rect 6472 16046 6500 16526
rect 6276 16040 6328 16046
rect 6276 15982 6328 15988
rect 6460 16040 6512 16046
rect 6460 15982 6512 15988
rect 6368 15904 6420 15910
rect 6368 15846 6420 15852
rect 6380 15434 6408 15846
rect 6472 15638 6500 15982
rect 6460 15632 6512 15638
rect 6460 15574 6512 15580
rect 6368 15428 6420 15434
rect 6368 15370 6420 15376
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6644 13932 6696 13938
rect 6644 13874 6696 13880
rect 6656 13802 6684 13874
rect 6748 13870 6776 14214
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 6644 13796 6696 13802
rect 6644 13738 6696 13744
rect 6656 13258 6684 13738
rect 6644 13252 6696 13258
rect 6644 13194 6696 13200
rect 6932 12850 6960 18634
rect 7024 17202 7052 18788
rect 7012 17196 7064 17202
rect 7012 17138 7064 17144
rect 7024 16726 7052 17138
rect 7012 16720 7064 16726
rect 7012 16662 7064 16668
rect 7024 14958 7052 16662
rect 7104 16652 7156 16658
rect 7104 16594 7156 16600
rect 7116 16114 7144 16594
rect 7104 16108 7156 16114
rect 7104 16050 7156 16056
rect 7208 16046 7236 19382
rect 7380 19372 7432 19378
rect 7380 19314 7432 19320
rect 7288 18828 7340 18834
rect 7288 18770 7340 18776
rect 7300 18222 7328 18770
rect 7392 18766 7420 19314
rect 7380 18760 7432 18766
rect 7380 18702 7432 18708
rect 7392 18290 7420 18702
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 7484 18222 7512 19910
rect 7656 19712 7708 19718
rect 7656 19654 7708 19660
rect 7668 19446 7696 19654
rect 7656 19440 7708 19446
rect 7656 19382 7708 19388
rect 8404 19310 8432 22066
rect 8576 22034 8628 22040
rect 8668 22092 8720 22098
rect 8668 22034 8720 22040
rect 9312 22092 9364 22098
rect 9496 22092 9548 22098
rect 9364 22052 9444 22080
rect 9312 22034 9364 22040
rect 8588 22001 8616 22034
rect 8574 21992 8630 22001
rect 8574 21927 8630 21936
rect 8576 21684 8628 21690
rect 8576 21626 8628 21632
rect 8588 21486 8616 21626
rect 8852 21616 8904 21622
rect 8852 21558 8904 21564
rect 8864 21486 8892 21558
rect 9220 21548 9272 21554
rect 9220 21490 9272 21496
rect 8576 21480 8628 21486
rect 8576 21422 8628 21428
rect 8852 21480 8904 21486
rect 8852 21422 8904 21428
rect 8944 21480 8996 21486
rect 8944 21422 8996 21428
rect 8576 21344 8628 21350
rect 8576 21286 8628 21292
rect 8668 21344 8720 21350
rect 8668 21286 8720 21292
rect 8484 21004 8536 21010
rect 8484 20946 8536 20952
rect 8392 19304 8444 19310
rect 8392 19246 8444 19252
rect 7564 19168 7616 19174
rect 7564 19110 7616 19116
rect 7576 18766 7604 19110
rect 7564 18760 7616 18766
rect 7564 18702 7616 18708
rect 8128 18686 8340 18714
rect 7288 18216 7340 18222
rect 7288 18158 7340 18164
rect 7472 18216 7524 18222
rect 7472 18158 7524 18164
rect 7380 18080 7432 18086
rect 7380 18022 7432 18028
rect 7748 18080 7800 18086
rect 7748 18022 7800 18028
rect 7196 16040 7248 16046
rect 7196 15982 7248 15988
rect 7208 15638 7236 15982
rect 7196 15632 7248 15638
rect 7196 15574 7248 15580
rect 7012 14952 7064 14958
rect 7012 14894 7064 14900
rect 7024 13394 7052 14894
rect 7208 14482 7236 15574
rect 7196 14476 7248 14482
rect 7196 14418 7248 14424
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7208 12306 7236 12786
rect 7392 12306 7420 18022
rect 7472 16992 7524 16998
rect 7472 16934 7524 16940
rect 7484 16658 7512 16934
rect 7760 16726 7788 18022
rect 8128 17202 8156 18686
rect 8312 18630 8340 18686
rect 8208 18624 8260 18630
rect 8208 18566 8260 18572
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 8116 17196 8168 17202
rect 8116 17138 8168 17144
rect 7748 16720 7800 16726
rect 7748 16662 7800 16668
rect 8116 16720 8168 16726
rect 8116 16662 8168 16668
rect 7472 16652 7524 16658
rect 7472 16594 7524 16600
rect 7748 16516 7800 16522
rect 7748 16458 7800 16464
rect 7760 16114 7788 16458
rect 7748 16108 7800 16114
rect 7748 16050 7800 16056
rect 8024 16108 8076 16114
rect 8024 16050 8076 16056
rect 7760 15570 7788 16050
rect 8036 15706 8064 16050
rect 8024 15700 8076 15706
rect 8024 15642 8076 15648
rect 7748 15564 7800 15570
rect 7748 15506 7800 15512
rect 8128 15502 8156 16662
rect 8220 16454 8248 18566
rect 8404 18222 8432 19246
rect 8496 18766 8524 20946
rect 8484 18760 8536 18766
rect 8484 18702 8536 18708
rect 8392 18216 8444 18222
rect 8392 18158 8444 18164
rect 8300 16720 8352 16726
rect 8300 16662 8352 16668
rect 8208 16448 8260 16454
rect 8208 16390 8260 16396
rect 8220 15570 8248 16390
rect 8312 16182 8340 16662
rect 8588 16538 8616 21286
rect 8680 21078 8708 21286
rect 8668 21072 8720 21078
rect 8668 21014 8720 21020
rect 8956 21010 8984 21422
rect 9036 21412 9088 21418
rect 9036 21354 9088 21360
rect 8944 21004 8996 21010
rect 8944 20946 8996 20952
rect 9048 20806 9076 21354
rect 9232 21010 9260 21490
rect 9416 21418 9444 22052
rect 9496 22034 9548 22040
rect 9508 21622 9536 22034
rect 9496 21616 9548 21622
rect 9496 21558 9548 21564
rect 9600 21554 9628 22918
rect 13820 22636 13872 22642
rect 13820 22578 13872 22584
rect 10600 22568 10652 22574
rect 10520 22528 10600 22556
rect 10416 22500 10468 22506
rect 10416 22442 10468 22448
rect 10324 22432 10376 22438
rect 10322 22400 10324 22409
rect 10376 22400 10378 22409
rect 10322 22335 10378 22344
rect 10232 21888 10284 21894
rect 10232 21830 10284 21836
rect 9772 21684 9824 21690
rect 9772 21626 9824 21632
rect 9588 21548 9640 21554
rect 9588 21490 9640 21496
rect 9312 21412 9364 21418
rect 9312 21354 9364 21360
rect 9404 21412 9456 21418
rect 9404 21354 9456 21360
rect 9324 21010 9352 21354
rect 9416 21321 9444 21354
rect 9402 21312 9458 21321
rect 9402 21247 9458 21256
rect 9784 21146 9812 21626
rect 10244 21554 10272 21830
rect 10232 21548 10284 21554
rect 10232 21490 10284 21496
rect 10336 21486 10364 22335
rect 10428 22098 10456 22442
rect 10520 22098 10548 22528
rect 10600 22510 10652 22516
rect 11796 22568 11848 22574
rect 11796 22510 11848 22516
rect 12532 22568 12584 22574
rect 12532 22510 12584 22516
rect 12808 22568 12860 22574
rect 12808 22510 12860 22516
rect 11704 22432 11756 22438
rect 11704 22374 11756 22380
rect 10416 22092 10468 22098
rect 10416 22034 10468 22040
rect 10508 22092 10560 22098
rect 10508 22034 10560 22040
rect 10784 22092 10836 22098
rect 10784 22034 10836 22040
rect 10428 21962 10456 22034
rect 10416 21956 10468 21962
rect 10416 21898 10468 21904
rect 10520 21690 10548 22034
rect 10692 22024 10744 22030
rect 10692 21966 10744 21972
rect 10508 21684 10560 21690
rect 10508 21626 10560 21632
rect 10704 21486 10732 21966
rect 10324 21480 10376 21486
rect 10324 21422 10376 21428
rect 10692 21480 10744 21486
rect 10692 21422 10744 21428
rect 10140 21344 10192 21350
rect 10140 21286 10192 21292
rect 10692 21344 10744 21350
rect 10796 21332 10824 22034
rect 11716 21962 11744 22374
rect 11808 22166 11836 22510
rect 12072 22500 12124 22506
rect 12072 22442 12124 22448
rect 12440 22500 12492 22506
rect 12440 22442 12492 22448
rect 11796 22160 11848 22166
rect 11796 22102 11848 22108
rect 11704 21956 11756 21962
rect 11704 21898 11756 21904
rect 11716 21865 11744 21898
rect 11702 21856 11758 21865
rect 11702 21791 11758 21800
rect 11716 21554 11744 21791
rect 11704 21548 11756 21554
rect 11704 21490 11756 21496
rect 11808 21486 11836 22102
rect 11796 21480 11848 21486
rect 11796 21422 11848 21428
rect 12084 21418 12112 22442
rect 12256 22432 12308 22438
rect 12256 22374 12308 22380
rect 12268 21554 12296 22374
rect 12452 21690 12480 22442
rect 12544 22234 12572 22510
rect 12716 22432 12768 22438
rect 12716 22374 12768 22380
rect 12532 22228 12584 22234
rect 12532 22170 12584 22176
rect 12440 21684 12492 21690
rect 12440 21626 12492 21632
rect 12532 21616 12584 21622
rect 12532 21558 12584 21564
rect 12256 21548 12308 21554
rect 12256 21490 12308 21496
rect 11336 21412 11388 21418
rect 11336 21354 11388 21360
rect 12072 21412 12124 21418
rect 12072 21354 12124 21360
rect 10744 21304 10824 21332
rect 11060 21344 11112 21350
rect 10692 21286 10744 21292
rect 11060 21286 11112 21292
rect 11152 21344 11204 21350
rect 11152 21286 11204 21292
rect 9772 21140 9824 21146
rect 9772 21082 9824 21088
rect 10152 21078 10180 21286
rect 10704 21146 10732 21286
rect 10692 21140 10744 21146
rect 10692 21082 10744 21088
rect 10140 21072 10192 21078
rect 10140 21014 10192 21020
rect 9128 21004 9180 21010
rect 9128 20946 9180 20952
rect 9220 21004 9272 21010
rect 9220 20946 9272 20952
rect 9312 21004 9364 21010
rect 9312 20946 9364 20952
rect 10048 21004 10100 21010
rect 10048 20946 10100 20952
rect 9036 20800 9088 20806
rect 9036 20742 9088 20748
rect 9048 20398 9076 20742
rect 9036 20392 9088 20398
rect 9036 20334 9088 20340
rect 8760 19916 8812 19922
rect 8760 19858 8812 19864
rect 8772 19310 8800 19858
rect 8760 19304 8812 19310
rect 8760 19246 8812 19252
rect 8772 18834 8800 19246
rect 9048 18902 9076 20334
rect 9140 19922 9168 20946
rect 9324 20788 9352 20946
rect 9404 20800 9456 20806
rect 9324 20760 9404 20788
rect 9404 20742 9456 20748
rect 10060 20602 10088 20946
rect 10692 20868 10744 20874
rect 10692 20810 10744 20816
rect 10048 20596 10100 20602
rect 10048 20538 10100 20544
rect 9588 20392 9640 20398
rect 9588 20334 9640 20340
rect 9128 19916 9180 19922
rect 9128 19858 9180 19864
rect 9496 19848 9548 19854
rect 9496 19790 9548 19796
rect 9508 19242 9536 19790
rect 9496 19236 9548 19242
rect 9496 19178 9548 19184
rect 9036 18896 9088 18902
rect 9036 18838 9088 18844
rect 9600 18834 9628 20334
rect 9864 19916 9916 19922
rect 9864 19858 9916 19864
rect 9876 19334 9904 19858
rect 9784 19306 9904 19334
rect 10704 19310 10732 20810
rect 10968 20596 11020 20602
rect 10968 20538 11020 20544
rect 10980 19310 11008 20538
rect 11072 19854 11100 21286
rect 11164 20806 11192 21286
rect 11152 20800 11204 20806
rect 11152 20742 11204 20748
rect 11244 19916 11296 19922
rect 11244 19858 11296 19864
rect 11060 19848 11112 19854
rect 11060 19790 11112 19796
rect 9784 19242 9812 19306
rect 10692 19304 10744 19310
rect 10692 19246 10744 19252
rect 10968 19304 11020 19310
rect 10968 19246 11020 19252
rect 9772 19236 9824 19242
rect 9772 19178 9824 19184
rect 10600 19236 10652 19242
rect 10600 19178 10652 19184
rect 10612 18834 10640 19178
rect 10704 18902 10732 19246
rect 10980 18902 11008 19246
rect 10692 18896 10744 18902
rect 10692 18838 10744 18844
rect 10968 18896 11020 18902
rect 10968 18838 11020 18844
rect 11072 18834 11100 19790
rect 8760 18828 8812 18834
rect 8760 18770 8812 18776
rect 9588 18828 9640 18834
rect 9588 18770 9640 18776
rect 10416 18828 10468 18834
rect 10416 18770 10468 18776
rect 10600 18828 10652 18834
rect 10600 18770 10652 18776
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 8772 18222 8800 18770
rect 9496 18692 9548 18698
rect 9496 18634 9548 18640
rect 8760 18216 8812 18222
rect 8760 18158 8812 18164
rect 9036 18148 9088 18154
rect 9036 18090 9088 18096
rect 8852 17128 8904 17134
rect 8852 17070 8904 17076
rect 8496 16510 8616 16538
rect 8864 16522 8892 17070
rect 8852 16516 8904 16522
rect 8300 16176 8352 16182
rect 8300 16118 8352 16124
rect 8312 15706 8340 16118
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8300 15700 8352 15706
rect 8300 15642 8352 15648
rect 8208 15564 8260 15570
rect 8208 15506 8260 15512
rect 8116 15496 8168 15502
rect 8116 15438 8168 15444
rect 8024 14476 8076 14482
rect 8024 14418 8076 14424
rect 8036 13870 8064 14418
rect 8404 14414 8432 15846
rect 8392 14408 8444 14414
rect 8392 14350 8444 14356
rect 8404 13870 8432 14350
rect 8024 13864 8076 13870
rect 8024 13806 8076 13812
rect 8392 13864 8444 13870
rect 8392 13806 8444 13812
rect 8208 13388 8260 13394
rect 8208 13330 8260 13336
rect 7932 12640 7984 12646
rect 7932 12582 7984 12588
rect 7196 12300 7248 12306
rect 7196 12242 7248 12248
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7208 11694 7236 12242
rect 7392 11694 7420 12242
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 7564 11824 7616 11830
rect 7564 11766 7616 11772
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7012 11620 7064 11626
rect 7012 11562 7064 11568
rect 6184 11348 6236 11354
rect 6184 11290 6236 11296
rect 7024 11286 7052 11562
rect 7012 11280 7064 11286
rect 7012 11222 7064 11228
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 5632 11008 5684 11014
rect 5632 10950 5684 10956
rect 5644 10606 5672 10950
rect 6748 10810 6776 11154
rect 6736 10804 6788 10810
rect 6736 10746 6788 10752
rect 5356 10600 5408 10606
rect 5356 10542 5408 10548
rect 5632 10600 5684 10606
rect 5632 10542 5684 10548
rect 5368 10130 5396 10542
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 4988 9648 5040 9654
rect 4988 9590 5040 9596
rect 5080 9648 5132 9654
rect 5080 9590 5132 9596
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 5000 8634 5028 8978
rect 5092 8838 5120 9590
rect 5460 9518 5488 10202
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 5460 8566 5488 9454
rect 5724 9376 5776 9382
rect 5724 9318 5776 9324
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 5736 8634 5764 9318
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5448 8560 5500 8566
rect 5448 8502 5500 8508
rect 4160 8356 4212 8362
rect 4160 8298 4212 8304
rect 4712 8356 4764 8362
rect 4712 8298 4764 8304
rect 4804 8356 4856 8362
rect 4804 8298 4856 8304
rect 5816 8356 5868 8362
rect 5816 8298 5868 8304
rect 4322 8188 4630 8197
rect 4322 8186 4328 8188
rect 4384 8186 4408 8188
rect 4464 8186 4488 8188
rect 4544 8186 4568 8188
rect 4624 8186 4630 8188
rect 4384 8134 4386 8186
rect 4566 8134 4568 8186
rect 4322 8132 4328 8134
rect 4384 8132 4408 8134
rect 4464 8132 4488 8134
rect 4544 8132 4568 8134
rect 4624 8132 4630 8134
rect 4322 8123 4630 8132
rect 4724 8090 4752 8298
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 4712 8084 4764 8090
rect 4712 8026 4764 8032
rect 3332 7948 3384 7954
rect 3332 7890 3384 7896
rect 3424 7948 3476 7954
rect 3424 7890 3476 7896
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 3068 7002 3096 7278
rect 3160 7262 3280 7290
rect 3056 6996 3108 7002
rect 3056 6938 3108 6944
rect 3252 6662 3280 7262
rect 3344 7206 3372 7890
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 3436 6934 3464 7890
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 3662 7644 3970 7653
rect 3662 7642 3668 7644
rect 3724 7642 3748 7644
rect 3804 7642 3828 7644
rect 3884 7642 3908 7644
rect 3964 7642 3970 7644
rect 3724 7590 3726 7642
rect 3906 7590 3908 7642
rect 3662 7588 3668 7590
rect 3724 7588 3748 7590
rect 3804 7588 3828 7590
rect 3884 7588 3908 7590
rect 3964 7588 3970 7590
rect 3662 7579 3970 7588
rect 3700 7268 3752 7274
rect 3700 7210 3752 7216
rect 3608 7200 3660 7206
rect 3608 7142 3660 7148
rect 3620 6934 3648 7142
rect 3712 7002 3740 7210
rect 3700 6996 3752 7002
rect 3700 6938 3752 6944
rect 3424 6928 3476 6934
rect 3424 6870 3476 6876
rect 3608 6928 3660 6934
rect 3608 6870 3660 6876
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 3436 5302 3464 6870
rect 3662 6556 3970 6565
rect 3662 6554 3668 6556
rect 3724 6554 3748 6556
rect 3804 6554 3828 6556
rect 3884 6554 3908 6556
rect 3964 6554 3970 6556
rect 3724 6502 3726 6554
rect 3906 6502 3908 6554
rect 3662 6500 3668 6502
rect 3724 6500 3748 6502
rect 3804 6500 3828 6502
rect 3884 6500 3908 6502
rect 3964 6500 3970 6502
rect 3662 6491 3970 6500
rect 4264 6390 4292 7686
rect 4724 7410 4752 8026
rect 4712 7404 4764 7410
rect 4712 7346 4764 7352
rect 4896 7336 4948 7342
rect 4896 7278 4948 7284
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4322 7100 4630 7109
rect 4322 7098 4328 7100
rect 4384 7098 4408 7100
rect 4464 7098 4488 7100
rect 4544 7098 4568 7100
rect 4624 7098 4630 7100
rect 4384 7046 4386 7098
rect 4566 7046 4568 7098
rect 4322 7044 4328 7046
rect 4384 7044 4408 7046
rect 4464 7044 4488 7046
rect 4544 7044 4568 7046
rect 4624 7044 4630 7046
rect 4322 7035 4630 7044
rect 4816 7018 4844 7142
rect 4724 6990 4844 7018
rect 4908 7002 4936 7278
rect 4896 6996 4948 7002
rect 4724 6458 4752 6990
rect 4896 6938 4948 6944
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4816 6458 4844 6802
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 4252 6384 4304 6390
rect 4252 6326 4304 6332
rect 3516 6112 3568 6118
rect 3516 6054 3568 6060
rect 3528 5370 3556 6054
rect 4264 5846 4292 6326
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 4322 6012 4630 6021
rect 4322 6010 4328 6012
rect 4384 6010 4408 6012
rect 4464 6010 4488 6012
rect 4544 6010 4568 6012
rect 4624 6010 4630 6012
rect 4384 5958 4386 6010
rect 4566 5958 4568 6010
rect 4322 5956 4328 5958
rect 4384 5956 4408 5958
rect 4464 5956 4488 5958
rect 4544 5956 4568 5958
rect 4624 5956 4630 5958
rect 4322 5947 4630 5956
rect 4252 5840 4304 5846
rect 4252 5782 4304 5788
rect 3662 5468 3970 5477
rect 3662 5466 3668 5468
rect 3724 5466 3748 5468
rect 3804 5466 3828 5468
rect 3884 5466 3908 5468
rect 3964 5466 3970 5468
rect 3724 5414 3726 5466
rect 3906 5414 3908 5466
rect 3662 5412 3668 5414
rect 3724 5412 3748 5414
rect 3804 5412 3828 5414
rect 3884 5412 3908 5414
rect 3964 5412 3970 5414
rect 3662 5403 3970 5412
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 3424 5296 3476 5302
rect 3424 5238 3476 5244
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 2884 4758 2912 5102
rect 3332 5092 3384 5098
rect 3332 5034 3384 5040
rect 3240 5024 3292 5030
rect 3240 4966 3292 4972
rect 2872 4752 2924 4758
rect 2872 4694 2924 4700
rect 3056 4684 3108 4690
rect 3056 4626 3108 4632
rect 3148 4684 3200 4690
rect 3148 4626 3200 4632
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 2320 4276 2372 4282
rect 2320 4218 2372 4224
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 1768 4072 1820 4078
rect 1768 4014 1820 4020
rect 2884 3602 2912 4218
rect 2964 4004 3016 4010
rect 2964 3946 3016 3952
rect 2976 3670 3004 3946
rect 2964 3664 3016 3670
rect 2964 3606 3016 3612
rect 3068 3602 3096 4626
rect 3160 4078 3188 4626
rect 3252 4146 3280 4966
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 3148 4072 3200 4078
rect 3148 4014 3200 4020
rect 3160 3670 3188 4014
rect 3344 3738 3372 5034
rect 3424 5024 3476 5030
rect 3700 5024 3752 5030
rect 3424 4966 3476 4972
rect 3528 4984 3700 5012
rect 3332 3732 3384 3738
rect 3332 3674 3384 3680
rect 3148 3664 3200 3670
rect 3148 3606 3200 3612
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 3056 3596 3108 3602
rect 3056 3538 3108 3544
rect 2884 3058 2912 3538
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 3160 2990 3188 3606
rect 3436 3194 3464 4966
rect 3528 3670 3556 4984
rect 3700 4966 3752 4972
rect 3896 4758 3924 5238
rect 5552 5166 5580 6054
rect 5644 5710 5672 6734
rect 5828 6390 5856 8298
rect 5920 7954 5948 8774
rect 6092 8560 6144 8566
rect 6092 8502 6144 8508
rect 5908 7948 5960 7954
rect 5908 7890 5960 7896
rect 6104 7750 6132 8502
rect 6288 8430 6316 9318
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 6380 8430 6408 8570
rect 6748 8430 6776 10746
rect 7024 10606 7052 11222
rect 7576 10606 7604 11766
rect 7852 10606 7880 12174
rect 7944 11694 7972 12582
rect 8220 12306 8248 13330
rect 8496 12730 8524 16510
rect 8852 16458 8904 16464
rect 8576 16448 8628 16454
rect 8576 16390 8628 16396
rect 8588 12850 8616 16390
rect 8864 16046 8892 16458
rect 9048 16250 9076 18090
rect 9508 17814 9536 18634
rect 9600 18358 9628 18770
rect 10048 18624 10100 18630
rect 10048 18566 10100 18572
rect 10060 18358 10088 18566
rect 9588 18352 9640 18358
rect 9588 18294 9640 18300
rect 10048 18352 10100 18358
rect 10048 18294 10100 18300
rect 9956 18284 10008 18290
rect 9956 18226 10008 18232
rect 9496 17808 9548 17814
rect 9496 17750 9548 17756
rect 9508 17678 9536 17750
rect 9588 17740 9640 17746
rect 9588 17682 9640 17688
rect 9496 17672 9548 17678
rect 9496 17614 9548 17620
rect 9600 17338 9628 17682
rect 9968 17678 9996 18226
rect 10060 18222 10088 18294
rect 10428 18222 10456 18770
rect 10048 18216 10100 18222
rect 10048 18158 10100 18164
rect 10416 18216 10468 18222
rect 10612 18204 10640 18770
rect 11256 18766 11284 19858
rect 11244 18760 11296 18766
rect 11244 18702 11296 18708
rect 10692 18216 10744 18222
rect 10612 18176 10692 18204
rect 10416 18158 10468 18164
rect 10692 18158 10744 18164
rect 11152 18216 11204 18222
rect 11152 18158 11204 18164
rect 9956 17672 10008 17678
rect 9956 17614 10008 17620
rect 9588 17332 9640 17338
rect 9588 17274 9640 17280
rect 9680 17332 9732 17338
rect 9680 17274 9732 17280
rect 9692 16794 9720 17274
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9692 16250 9720 16526
rect 9036 16244 9088 16250
rect 9036 16186 9088 16192
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9048 16046 9076 16186
rect 8668 16040 8720 16046
rect 8668 15982 8720 15988
rect 8852 16040 8904 16046
rect 8852 15982 8904 15988
rect 9036 16040 9088 16046
rect 9036 15982 9088 15988
rect 8680 15434 8708 15982
rect 8668 15428 8720 15434
rect 8668 15370 8720 15376
rect 8760 15360 8812 15366
rect 8760 15302 8812 15308
rect 8668 13728 8720 13734
rect 8668 13670 8720 13676
rect 8576 12844 8628 12850
rect 8576 12786 8628 12792
rect 8404 12714 8524 12730
rect 8392 12708 8524 12714
rect 8444 12702 8524 12708
rect 8392 12650 8444 12656
rect 8588 12374 8616 12786
rect 8680 12782 8708 13670
rect 8772 12986 8800 15302
rect 10060 14550 10088 18158
rect 11060 18148 11112 18154
rect 11060 18090 11112 18096
rect 11072 16726 11100 18090
rect 11164 17882 11192 18158
rect 11152 17876 11204 17882
rect 11152 17818 11204 17824
rect 11060 16720 11112 16726
rect 11060 16662 11112 16668
rect 10968 16584 11020 16590
rect 10968 16526 11020 16532
rect 10980 16250 11008 16526
rect 10968 16244 11020 16250
rect 10968 16186 11020 16192
rect 10968 16040 11020 16046
rect 10968 15982 11020 15988
rect 10980 15502 11008 15982
rect 11072 15978 11100 16662
rect 11060 15972 11112 15978
rect 11060 15914 11112 15920
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 10980 15094 11008 15438
rect 10968 15088 11020 15094
rect 10968 15030 11020 15036
rect 11072 14958 11100 15914
rect 11348 15570 11376 21354
rect 12268 21010 12296 21490
rect 12544 21350 12572 21558
rect 12728 21554 12756 22374
rect 12820 22098 12848 22510
rect 12900 22500 12952 22506
rect 12900 22442 12952 22448
rect 12912 22098 12940 22442
rect 13360 22228 13412 22234
rect 13360 22170 13412 22176
rect 13372 22098 13400 22170
rect 13728 22160 13780 22166
rect 13648 22120 13728 22148
rect 12808 22092 12860 22098
rect 12808 22034 12860 22040
rect 12900 22092 12952 22098
rect 12900 22034 12952 22040
rect 13360 22092 13412 22098
rect 13360 22034 13412 22040
rect 13268 22024 13320 22030
rect 13268 21966 13320 21972
rect 12900 21684 12952 21690
rect 12900 21626 12952 21632
rect 12716 21548 12768 21554
rect 12716 21490 12768 21496
rect 12808 21480 12860 21486
rect 12808 21422 12860 21428
rect 12532 21344 12584 21350
rect 12532 21286 12584 21292
rect 12820 21010 12848 21422
rect 12912 21418 12940 21626
rect 13280 21486 13308 21966
rect 13648 21690 13676 22120
rect 13728 22102 13780 22108
rect 13832 22030 13860 22578
rect 13924 22234 13952 23054
rect 14096 22976 14148 22982
rect 14096 22918 14148 22924
rect 14004 22772 14056 22778
rect 14004 22714 14056 22720
rect 13912 22228 13964 22234
rect 13912 22170 13964 22176
rect 14016 22098 14044 22714
rect 14108 22574 14136 22918
rect 14096 22568 14148 22574
rect 14096 22510 14148 22516
rect 15212 22506 15240 23054
rect 15292 22772 15344 22778
rect 15292 22714 15344 22720
rect 15304 22574 15332 22714
rect 15292 22568 15344 22574
rect 15292 22510 15344 22516
rect 14188 22500 14240 22506
rect 14188 22442 14240 22448
rect 15200 22500 15252 22506
rect 15200 22442 15252 22448
rect 14096 22228 14148 22234
rect 14096 22170 14148 22176
rect 14004 22092 14056 22098
rect 14004 22034 14056 22040
rect 13820 22024 13872 22030
rect 13820 21966 13872 21972
rect 13728 21888 13780 21894
rect 13728 21830 13780 21836
rect 13636 21684 13688 21690
rect 13636 21626 13688 21632
rect 13740 21554 13768 21830
rect 14108 21622 14136 22170
rect 14200 21894 14228 22442
rect 14832 22432 14884 22438
rect 14646 22400 14702 22409
rect 14832 22374 14884 22380
rect 15016 22432 15068 22438
rect 15016 22374 15068 22380
rect 14646 22335 14702 22344
rect 14660 21962 14688 22335
rect 14740 22160 14792 22166
rect 14740 22102 14792 22108
rect 14648 21956 14700 21962
rect 14648 21898 14700 21904
rect 14188 21888 14240 21894
rect 14188 21830 14240 21836
rect 14096 21616 14148 21622
rect 14096 21558 14148 21564
rect 13728 21548 13780 21554
rect 13728 21490 13780 21496
rect 13268 21480 13320 21486
rect 13268 21422 13320 21428
rect 12900 21412 12952 21418
rect 12900 21354 12952 21360
rect 13544 21412 13596 21418
rect 13544 21354 13596 21360
rect 13084 21344 13136 21350
rect 13084 21286 13136 21292
rect 13360 21344 13412 21350
rect 13360 21286 13412 21292
rect 13096 21010 13124 21286
rect 12256 21004 12308 21010
rect 12256 20946 12308 20952
rect 12808 21004 12860 21010
rect 12808 20946 12860 20952
rect 13084 21004 13136 21010
rect 13084 20946 13136 20952
rect 12808 20800 12860 20806
rect 12808 20742 12860 20748
rect 11520 19712 11572 19718
rect 11520 19654 11572 19660
rect 11532 19378 11560 19654
rect 11520 19372 11572 19378
rect 11520 19314 11572 19320
rect 12164 19372 12216 19378
rect 12164 19314 12216 19320
rect 12176 18834 12204 19314
rect 12256 18964 12308 18970
rect 12256 18906 12308 18912
rect 12164 18828 12216 18834
rect 12164 18770 12216 18776
rect 12268 18154 12296 18906
rect 12716 18828 12768 18834
rect 12716 18770 12768 18776
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12440 18352 12492 18358
rect 12440 18294 12492 18300
rect 12256 18148 12308 18154
rect 12256 18090 12308 18096
rect 12164 18080 12216 18086
rect 12164 18022 12216 18028
rect 11520 16992 11572 16998
rect 11520 16934 11572 16940
rect 11532 16794 11560 16934
rect 11520 16788 11572 16794
rect 11520 16730 11572 16736
rect 12176 16658 12204 18022
rect 12452 17746 12480 18294
rect 12544 18222 12572 18702
rect 12624 18624 12676 18630
rect 12624 18566 12676 18572
rect 12636 18426 12664 18566
rect 12624 18420 12676 18426
rect 12624 18362 12676 18368
rect 12728 18290 12756 18770
rect 12716 18284 12768 18290
rect 12716 18226 12768 18232
rect 12532 18216 12584 18222
rect 12532 18158 12584 18164
rect 12440 17740 12492 17746
rect 12440 17682 12492 17688
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 12164 16652 12216 16658
rect 12164 16594 12216 16600
rect 12360 16590 12388 16730
rect 12348 16584 12400 16590
rect 12348 16526 12400 16532
rect 12624 16176 12676 16182
rect 12624 16118 12676 16124
rect 11612 15972 11664 15978
rect 11612 15914 11664 15920
rect 11624 15706 11652 15914
rect 11612 15700 11664 15706
rect 11612 15642 11664 15648
rect 11336 15564 11388 15570
rect 11336 15506 11388 15512
rect 11244 15496 11296 15502
rect 11244 15438 11296 15444
rect 11256 15162 11284 15438
rect 11244 15156 11296 15162
rect 11244 15098 11296 15104
rect 12636 14958 12664 16118
rect 12820 16046 12848 20742
rect 13176 19372 13228 19378
rect 13176 19314 13228 19320
rect 12992 19304 13044 19310
rect 12992 19246 13044 19252
rect 13004 18834 13032 19246
rect 12992 18828 13044 18834
rect 12992 18770 13044 18776
rect 12900 18624 12952 18630
rect 12900 18566 12952 18572
rect 12912 18306 12940 18566
rect 13084 18352 13136 18358
rect 12912 18300 13084 18306
rect 12912 18294 13136 18300
rect 12912 18278 13124 18294
rect 12912 17542 12940 18278
rect 13188 17746 13216 19314
rect 13268 19304 13320 19310
rect 13372 19292 13400 21286
rect 13320 19264 13400 19292
rect 13268 19246 13320 19252
rect 13372 18834 13400 19264
rect 13360 18828 13412 18834
rect 13360 18770 13412 18776
rect 13268 18760 13320 18766
rect 13268 18702 13320 18708
rect 13280 18290 13308 18702
rect 13268 18284 13320 18290
rect 13268 18226 13320 18232
rect 13452 18148 13504 18154
rect 13452 18090 13504 18096
rect 13464 17814 13492 18090
rect 13452 17808 13504 17814
rect 13452 17750 13504 17756
rect 13176 17740 13228 17746
rect 13176 17682 13228 17688
rect 12900 17536 12952 17542
rect 12900 17478 12952 17484
rect 13188 17134 13216 17682
rect 13556 17354 13584 21354
rect 14200 21146 14228 21830
rect 14752 21690 14780 22102
rect 14740 21684 14792 21690
rect 14740 21626 14792 21632
rect 14844 21486 14872 22374
rect 15028 22234 15056 22374
rect 15016 22228 15068 22234
rect 15016 22170 15068 22176
rect 15016 21956 15068 21962
rect 15016 21898 15068 21904
rect 14832 21480 14884 21486
rect 14832 21422 14884 21428
rect 14740 21412 14792 21418
rect 14740 21354 14792 21360
rect 14188 21140 14240 21146
rect 14188 21082 14240 21088
rect 14752 21010 14780 21354
rect 14844 21078 14872 21422
rect 15028 21146 15056 21898
rect 15108 21480 15160 21486
rect 15108 21422 15160 21428
rect 15016 21140 15068 21146
rect 15016 21082 15068 21088
rect 14832 21072 14884 21078
rect 14832 21014 14884 21020
rect 14740 21004 14792 21010
rect 14740 20946 14792 20952
rect 14188 20936 14240 20942
rect 14188 20878 14240 20884
rect 13912 18692 13964 18698
rect 13912 18634 13964 18640
rect 13924 18086 13952 18634
rect 13912 18080 13964 18086
rect 13912 18022 13964 18028
rect 14004 18080 14056 18086
rect 14004 18022 14056 18028
rect 13924 17814 13952 18022
rect 13912 17808 13964 17814
rect 13912 17750 13964 17756
rect 14016 17746 14044 18022
rect 14004 17740 14056 17746
rect 14004 17682 14056 17688
rect 13912 17672 13964 17678
rect 13464 17326 13584 17354
rect 13740 17620 13912 17626
rect 13740 17614 13964 17620
rect 13740 17598 13952 17614
rect 13176 17128 13228 17134
rect 13176 17070 13228 17076
rect 13464 16046 13492 17326
rect 13544 17196 13596 17202
rect 13544 17138 13596 17144
rect 13556 16250 13584 17138
rect 13740 17134 13768 17598
rect 14004 17536 14056 17542
rect 14004 17478 14056 17484
rect 13728 17128 13780 17134
rect 13728 17070 13780 17076
rect 13636 17060 13688 17066
rect 13636 17002 13688 17008
rect 13648 16726 13676 17002
rect 14016 16726 14044 17478
rect 14096 17196 14148 17202
rect 14096 17138 14148 17144
rect 13636 16720 13688 16726
rect 13636 16662 13688 16668
rect 14004 16720 14056 16726
rect 14004 16662 14056 16668
rect 13728 16652 13780 16658
rect 13728 16594 13780 16600
rect 13912 16652 13964 16658
rect 13912 16594 13964 16600
rect 13544 16244 13596 16250
rect 13544 16186 13596 16192
rect 13740 16046 13768 16594
rect 13924 16046 13952 16594
rect 14016 16114 14044 16662
rect 14004 16108 14056 16114
rect 14004 16050 14056 16056
rect 12808 16040 12860 16046
rect 12808 15982 12860 15988
rect 13268 16040 13320 16046
rect 13452 16040 13504 16046
rect 13268 15982 13320 15988
rect 13372 16000 13452 16028
rect 13176 15904 13228 15910
rect 13176 15846 13228 15852
rect 12900 15428 12952 15434
rect 12900 15370 12952 15376
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 12624 14952 12676 14958
rect 12624 14894 12676 14900
rect 10048 14544 10100 14550
rect 10048 14486 10100 14492
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 8944 14272 8996 14278
rect 8944 14214 8996 14220
rect 8852 14000 8904 14006
rect 8852 13942 8904 13948
rect 8864 13802 8892 13942
rect 8956 13938 8984 14214
rect 8944 13932 8996 13938
rect 8944 13874 8996 13880
rect 9048 13870 9076 14418
rect 9680 14340 9732 14346
rect 9680 14282 9732 14288
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 9036 13864 9088 13870
rect 9036 13806 9088 13812
rect 8852 13796 8904 13802
rect 8852 13738 8904 13744
rect 9508 13462 9536 14010
rect 9496 13456 9548 13462
rect 9496 13398 9548 13404
rect 9692 13326 9720 14282
rect 11072 13870 11100 14894
rect 11520 14816 11572 14822
rect 11520 14758 11572 14764
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 11244 14068 11296 14074
rect 11244 14010 11296 14016
rect 11256 13870 11284 14010
rect 11532 13870 11560 14758
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 11244 13864 11296 13870
rect 11244 13806 11296 13812
rect 11520 13864 11572 13870
rect 11520 13806 11572 13812
rect 12348 13796 12400 13802
rect 12348 13738 12400 13744
rect 10232 13728 10284 13734
rect 10232 13670 10284 13676
rect 10244 13394 10272 13670
rect 12360 13394 12388 13738
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 12728 13394 12756 13670
rect 12820 13394 12848 14758
rect 12912 13870 12940 15370
rect 12900 13864 12952 13870
rect 12900 13806 12952 13812
rect 12912 13530 12940 13806
rect 12900 13524 12952 13530
rect 12900 13466 12952 13472
rect 12912 13394 12940 13466
rect 13188 13394 13216 15846
rect 13280 15570 13308 15982
rect 13268 15564 13320 15570
rect 13268 15506 13320 15512
rect 13372 15502 13400 16000
rect 13452 15982 13504 15988
rect 13728 16040 13780 16046
rect 13728 15982 13780 15988
rect 13912 16040 13964 16046
rect 13912 15982 13964 15988
rect 13740 15910 13768 15982
rect 13452 15904 13504 15910
rect 13452 15846 13504 15852
rect 13728 15904 13780 15910
rect 13728 15846 13780 15852
rect 13464 15570 13492 15846
rect 13740 15706 13768 15846
rect 13728 15700 13780 15706
rect 13728 15642 13780 15648
rect 13452 15564 13504 15570
rect 13452 15506 13504 15512
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 13360 15496 13412 15502
rect 13360 15438 13412 15444
rect 13832 15162 13860 15506
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 13280 13394 13308 13874
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13648 13462 13676 13806
rect 13832 13530 13860 15098
rect 13924 14074 13952 15982
rect 13912 14068 13964 14074
rect 13912 14010 13964 14016
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13636 13456 13688 13462
rect 13636 13398 13688 13404
rect 10232 13388 10284 13394
rect 10232 13330 10284 13336
rect 12348 13388 12400 13394
rect 12348 13330 12400 13336
rect 12716 13388 12768 13394
rect 12716 13330 12768 13336
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12900 13388 12952 13394
rect 12900 13330 12952 13336
rect 13176 13388 13228 13394
rect 13176 13330 13228 13336
rect 13268 13388 13320 13394
rect 13268 13330 13320 13336
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9692 13190 9720 13262
rect 12360 13258 12388 13330
rect 9956 13252 10008 13258
rect 9956 13194 10008 13200
rect 12348 13252 12400 13258
rect 12348 13194 12400 13200
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 8576 12368 8628 12374
rect 8576 12310 8628 12316
rect 8772 12306 8800 12922
rect 9416 12782 9444 12922
rect 9680 12912 9732 12918
rect 9680 12854 9732 12860
rect 8852 12776 8904 12782
rect 8852 12718 8904 12724
rect 9404 12776 9456 12782
rect 9404 12718 9456 12724
rect 8864 12374 8892 12718
rect 9404 12640 9456 12646
rect 9404 12582 9456 12588
rect 9416 12442 9444 12582
rect 9404 12436 9456 12442
rect 9404 12378 9456 12384
rect 8852 12368 8904 12374
rect 8852 12310 8904 12316
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 8760 12300 8812 12306
rect 8760 12242 8812 12248
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 8404 11694 8432 12038
rect 9324 11694 9352 12038
rect 9416 11694 9444 12378
rect 9692 12374 9720 12854
rect 9680 12368 9732 12374
rect 9680 12310 9732 12316
rect 9692 12102 9720 12310
rect 9968 12306 9996 13194
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 10508 13184 10560 13190
rect 10508 13126 10560 13132
rect 10428 12850 10456 13126
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 10520 12306 10548 13126
rect 12256 12844 12308 12850
rect 12256 12786 12308 12792
rect 11888 12776 11940 12782
rect 11888 12718 11940 12724
rect 10692 12708 10744 12714
rect 10692 12650 10744 12656
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 10232 12300 10284 12306
rect 10232 12242 10284 12248
rect 10508 12300 10560 12306
rect 10508 12242 10560 12248
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 7932 11688 7984 11694
rect 7932 11630 7984 11636
rect 8392 11688 8444 11694
rect 8392 11630 8444 11636
rect 9312 11688 9364 11694
rect 9312 11630 9364 11636
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 8024 11552 8076 11558
rect 8024 11494 8076 11500
rect 8760 11552 8812 11558
rect 8760 11494 8812 11500
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 8036 11218 8064 11494
rect 8772 11218 8800 11494
rect 8024 11212 8076 11218
rect 8024 11154 8076 11160
rect 8760 11212 8812 11218
rect 8760 11154 8812 11160
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 8128 10810 8156 10950
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 8772 10606 8800 11154
rect 9140 10606 9168 11494
rect 7012 10600 7064 10606
rect 7012 10542 7064 10548
rect 7564 10600 7616 10606
rect 7564 10542 7616 10548
rect 7840 10600 7892 10606
rect 7840 10542 7892 10548
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 7288 10532 7340 10538
rect 7288 10474 7340 10480
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 7024 10198 7052 10406
rect 7300 10266 7328 10474
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 7012 10192 7064 10198
rect 7012 10134 7064 10140
rect 7760 8634 7788 10202
rect 7852 10130 7880 10542
rect 8116 10532 8168 10538
rect 8116 10474 8168 10480
rect 9404 10532 9456 10538
rect 9404 10474 9456 10480
rect 8128 10266 8156 10474
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 7840 10124 7892 10130
rect 7840 10066 7892 10072
rect 8864 9586 8892 10406
rect 9416 10062 9444 10474
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 8852 9580 8904 9586
rect 8852 9522 8904 9528
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 8404 9110 8432 9318
rect 8772 9178 8800 9318
rect 8760 9172 8812 9178
rect 8760 9114 8812 9120
rect 8392 9104 8444 9110
rect 8392 9046 8444 9052
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 8772 8498 8800 9114
rect 9416 9042 9444 9998
rect 8852 9036 8904 9042
rect 8852 8978 8904 8984
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 6276 8424 6328 8430
rect 6276 8366 6328 8372
rect 6368 8424 6420 8430
rect 6368 8366 6420 8372
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6184 8288 6236 8294
rect 6184 8230 6236 8236
rect 6196 7954 6224 8230
rect 6184 7948 6236 7954
rect 6184 7890 6236 7896
rect 6380 7886 6408 8366
rect 6748 7954 6776 8366
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 6736 7948 6788 7954
rect 6736 7890 6788 7896
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 6092 7744 6144 7750
rect 6092 7686 6144 7692
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6932 7410 6960 7686
rect 7392 7546 7420 7822
rect 7380 7540 7432 7546
rect 7380 7482 7432 7488
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 7196 7336 7248 7342
rect 7196 7278 7248 7284
rect 7760 7290 7788 8230
rect 8220 7886 8248 8230
rect 8772 7954 8800 8434
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 8760 7948 8812 7954
rect 8760 7890 8812 7896
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 7944 7546 7972 7686
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 8220 7478 8248 7822
rect 8404 7546 8432 7890
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8208 7472 8260 7478
rect 8208 7414 8260 7420
rect 8208 7336 8260 7342
rect 7760 7284 8208 7290
rect 7760 7278 8260 7284
rect 5816 6384 5868 6390
rect 5816 6326 5868 6332
rect 6828 6384 6880 6390
rect 6828 6326 6880 6332
rect 5828 6254 5856 6326
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 5816 6248 5868 6254
rect 5816 6190 5868 6196
rect 6552 6248 6604 6254
rect 6552 6190 6604 6196
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5736 5914 5764 6054
rect 5724 5908 5776 5914
rect 5724 5850 5776 5856
rect 5828 5846 5856 6190
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6460 6112 6512 6118
rect 6460 6054 6512 6060
rect 5816 5840 5868 5846
rect 5816 5782 5868 5788
rect 6380 5778 6408 6054
rect 6368 5772 6420 5778
rect 6368 5714 6420 5720
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 5644 5370 5672 5646
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 4322 4924 4630 4933
rect 4322 4922 4328 4924
rect 4384 4922 4408 4924
rect 4464 4922 4488 4924
rect 4544 4922 4568 4924
rect 4624 4922 4630 4924
rect 4384 4870 4386 4922
rect 4566 4870 4568 4922
rect 4322 4868 4328 4870
rect 4384 4868 4408 4870
rect 4464 4868 4488 4870
rect 4544 4868 4568 4870
rect 4624 4868 4630 4870
rect 4322 4859 4630 4868
rect 5644 4842 5672 5306
rect 6472 5098 6500 6054
rect 6460 5092 6512 5098
rect 6460 5034 6512 5040
rect 4068 4820 4120 4826
rect 5644 4814 5764 4842
rect 6564 4826 6592 6190
rect 6748 6118 6776 6258
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6748 5846 6776 6054
rect 6736 5840 6788 5846
rect 6736 5782 6788 5788
rect 6840 5370 6868 6326
rect 7208 6254 7236 7278
rect 7656 7268 7708 7274
rect 7760 7262 8248 7278
rect 7656 7210 7708 7216
rect 7668 6254 7696 7210
rect 8220 7206 8248 7262
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7656 6248 7708 6254
rect 7656 6190 7708 6196
rect 7208 5914 7236 6190
rect 7392 6118 7420 6190
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 4068 4762 4120 4768
rect 3884 4752 3936 4758
rect 3884 4694 3936 4700
rect 3662 4380 3970 4389
rect 3662 4378 3668 4380
rect 3724 4378 3748 4380
rect 3804 4378 3828 4380
rect 3884 4378 3908 4380
rect 3964 4378 3970 4380
rect 3724 4326 3726 4378
rect 3906 4326 3908 4378
rect 3662 4324 3668 4326
rect 3724 4324 3748 4326
rect 3804 4324 3828 4326
rect 3884 4324 3908 4326
rect 3964 4324 3970 4326
rect 3662 4315 3970 4324
rect 4080 4214 4108 4762
rect 5736 4758 5764 4814
rect 6552 4820 6604 4826
rect 6552 4762 6604 4768
rect 6840 4758 6868 5306
rect 7208 5166 7236 5850
rect 7196 5160 7248 5166
rect 7196 5102 7248 5108
rect 4712 4752 4764 4758
rect 4712 4694 4764 4700
rect 5632 4752 5684 4758
rect 5632 4694 5684 4700
rect 5724 4752 5776 4758
rect 5724 4694 5776 4700
rect 6828 4752 6880 4758
rect 6828 4694 6880 4700
rect 4160 4684 4212 4690
rect 4160 4626 4212 4632
rect 4068 4208 4120 4214
rect 4068 4150 4120 4156
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 3516 3664 3568 3670
rect 3516 3606 3568 3612
rect 4080 3602 4108 4014
rect 4172 4010 4200 4626
rect 4436 4548 4488 4554
rect 4436 4490 4488 4496
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 4356 4078 4384 4422
rect 4448 4282 4476 4490
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 4344 4072 4396 4078
rect 4344 4014 4396 4020
rect 4160 4004 4212 4010
rect 4160 3946 4212 3952
rect 4172 3670 4200 3946
rect 4322 3836 4630 3845
rect 4322 3834 4328 3836
rect 4384 3834 4408 3836
rect 4464 3834 4488 3836
rect 4544 3834 4568 3836
rect 4624 3834 4630 3836
rect 4384 3782 4386 3834
rect 4566 3782 4568 3834
rect 4322 3780 4328 3782
rect 4384 3780 4408 3782
rect 4464 3780 4488 3782
rect 4544 3780 4568 3782
rect 4624 3780 4630 3782
rect 4322 3771 4630 3780
rect 4724 3738 4752 4694
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 4816 4078 4844 4218
rect 5644 4146 5672 4694
rect 7208 4486 7236 5102
rect 7392 5030 7420 6054
rect 7668 5914 7696 6190
rect 8024 6112 8076 6118
rect 8024 6054 8076 6060
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7668 5250 7696 5850
rect 8036 5370 8064 6054
rect 8864 5778 8892 8978
rect 9496 7812 9548 7818
rect 9496 7754 9548 7760
rect 9508 6798 9536 7754
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 9784 6934 9812 7686
rect 9772 6928 9824 6934
rect 9772 6870 9824 6876
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9404 5908 9456 5914
rect 9404 5850 9456 5856
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 8852 5772 8904 5778
rect 8852 5714 8904 5720
rect 8312 5370 8340 5714
rect 8760 5568 8812 5574
rect 8760 5510 8812 5516
rect 8772 5370 8800 5510
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 8864 5250 8892 5714
rect 7576 5222 7696 5250
rect 8772 5234 8892 5250
rect 8772 5228 8904 5234
rect 8772 5222 8852 5228
rect 7576 5166 7604 5222
rect 7564 5160 7616 5166
rect 7564 5102 7616 5108
rect 8024 5092 8076 5098
rect 8024 5034 8076 5040
rect 8576 5092 8628 5098
rect 8576 5034 8628 5040
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7392 4622 7420 4966
rect 8036 4826 8064 5034
rect 8588 4826 8616 5034
rect 8024 4820 8076 4826
rect 8024 4762 8076 4768
rect 8576 4820 8628 4826
rect 8576 4762 8628 4768
rect 8772 4690 8800 5222
rect 8852 5170 8904 5176
rect 9416 5166 9444 5850
rect 9876 5778 9904 11698
rect 9968 11694 9996 12242
rect 10244 11898 10272 12242
rect 10704 12170 10732 12650
rect 11900 12646 11928 12718
rect 11704 12640 11756 12646
rect 11704 12582 11756 12588
rect 11888 12640 11940 12646
rect 11888 12582 11940 12588
rect 10692 12164 10744 12170
rect 10692 12106 10744 12112
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 10520 11762 10548 12038
rect 10704 11762 10732 12106
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 10692 11620 10744 11626
rect 10692 11562 10744 11568
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10428 10606 10456 11494
rect 10508 11212 10560 11218
rect 10508 11154 10560 11160
rect 10520 10810 10548 11154
rect 10704 11150 10732 11562
rect 10888 11354 10916 11630
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 11716 11218 11744 12582
rect 12268 11354 12296 12786
rect 12360 12306 12388 13194
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12532 12980 12584 12986
rect 12532 12922 12584 12928
rect 12452 12782 12480 12922
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12452 12442 12480 12582
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 12256 11348 12308 11354
rect 12256 11290 12308 11296
rect 12452 11218 12480 12378
rect 12544 12306 12572 12922
rect 12728 12782 12756 13330
rect 12820 12850 12848 13330
rect 13280 12986 13308 13330
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 12808 12844 12860 12850
rect 12808 12786 12860 12792
rect 12716 12776 12768 12782
rect 12716 12718 12768 12724
rect 13268 12640 13320 12646
rect 13268 12582 13320 12588
rect 13280 12306 13308 12582
rect 13372 12306 13400 13126
rect 13452 12844 13504 12850
rect 13452 12786 13504 12792
rect 13464 12306 13492 12786
rect 13832 12782 13860 13126
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 12532 12300 12584 12306
rect 12532 12242 12584 12248
rect 13268 12300 13320 12306
rect 13268 12242 13320 12248
rect 13360 12300 13412 12306
rect 13360 12242 13412 12248
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 13544 12232 13596 12238
rect 13544 12174 13596 12180
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 13096 11694 13124 12038
rect 13084 11688 13136 11694
rect 13084 11630 13136 11636
rect 13556 11354 13584 12174
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 12440 11212 12492 11218
rect 12440 11154 12492 11160
rect 10692 11144 10744 11150
rect 10692 11086 10744 11092
rect 10508 10804 10560 10810
rect 10508 10746 10560 10752
rect 10416 10600 10468 10606
rect 10416 10542 10468 10548
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 10520 9586 10548 10406
rect 10704 9586 10732 11086
rect 11256 10810 11284 11154
rect 13648 11150 13676 11494
rect 12900 11144 12952 11150
rect 12900 11086 12952 11092
rect 13636 11144 13688 11150
rect 13636 11086 13688 11092
rect 11612 11008 11664 11014
rect 11612 10950 11664 10956
rect 10968 10804 11020 10810
rect 10968 10746 11020 10752
rect 11244 10804 11296 10810
rect 11244 10746 11296 10752
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10060 9110 10088 9318
rect 10796 9178 10824 9318
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 10048 9104 10100 9110
rect 10048 9046 10100 9052
rect 10796 8498 10824 9114
rect 10980 8838 11008 10746
rect 11256 8974 11284 10746
rect 11624 10606 11652 10950
rect 11612 10600 11664 10606
rect 11612 10542 11664 10548
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12728 9722 12756 9862
rect 12716 9716 12768 9722
rect 12716 9658 12768 9664
rect 12912 9518 12940 11086
rect 14108 10674 14136 17138
rect 14200 14958 14228 20878
rect 14752 20330 14780 20946
rect 15120 20398 15148 21422
rect 15108 20392 15160 20398
rect 15108 20334 15160 20340
rect 14740 20324 14792 20330
rect 14740 20266 14792 20272
rect 15212 19242 15240 22442
rect 15292 22432 15344 22438
rect 15292 22374 15344 22380
rect 15304 22030 15332 22374
rect 15488 22166 15516 23054
rect 16672 22976 16724 22982
rect 16672 22918 16724 22924
rect 16684 22506 16712 22918
rect 17972 22778 18000 23122
rect 18420 23112 18472 23118
rect 18420 23054 18472 23060
rect 18328 22976 18380 22982
rect 18328 22918 18380 22924
rect 17960 22772 18012 22778
rect 17960 22714 18012 22720
rect 16856 22568 16908 22574
rect 16856 22510 16908 22516
rect 15660 22500 15712 22506
rect 15660 22442 15712 22448
rect 16672 22500 16724 22506
rect 16672 22442 16724 22448
rect 15672 22234 15700 22442
rect 15660 22228 15712 22234
rect 15660 22170 15712 22176
rect 15476 22160 15528 22166
rect 15476 22102 15528 22108
rect 15672 22098 15700 22170
rect 16868 22098 16896 22510
rect 16948 22228 17000 22234
rect 16948 22170 17000 22176
rect 15660 22092 15712 22098
rect 15660 22034 15712 22040
rect 16856 22092 16908 22098
rect 16856 22034 16908 22040
rect 15292 22024 15344 22030
rect 15292 21966 15344 21972
rect 16672 22024 16724 22030
rect 16672 21966 16724 21972
rect 15304 21418 15332 21966
rect 16304 21888 16356 21894
rect 16304 21830 16356 21836
rect 15568 21684 15620 21690
rect 15568 21626 15620 21632
rect 15580 21554 15608 21626
rect 15568 21548 15620 21554
rect 15568 21490 15620 21496
rect 15292 21412 15344 21418
rect 15292 21354 15344 21360
rect 16028 21412 16080 21418
rect 16028 21354 16080 21360
rect 15568 21344 15620 21350
rect 15568 21286 15620 21292
rect 15936 21344 15988 21350
rect 15936 21286 15988 21292
rect 15580 21146 15608 21286
rect 15568 21140 15620 21146
rect 15568 21082 15620 21088
rect 15580 21010 15608 21082
rect 15948 21010 15976 21286
rect 16040 21078 16068 21354
rect 16028 21072 16080 21078
rect 16028 21014 16080 21020
rect 15568 21004 15620 21010
rect 15568 20946 15620 20952
rect 15936 21004 15988 21010
rect 15936 20946 15988 20952
rect 16316 20874 16344 21830
rect 16304 20868 16356 20874
rect 16304 20810 16356 20816
rect 16212 20800 16264 20806
rect 16212 20742 16264 20748
rect 16224 19310 16252 20742
rect 16684 20398 16712 21966
rect 16764 21684 16816 21690
rect 16764 21626 16816 21632
rect 16776 21010 16804 21626
rect 16960 21486 16988 22170
rect 17972 22098 18000 22714
rect 18340 22642 18368 22918
rect 18328 22636 18380 22642
rect 18328 22578 18380 22584
rect 18432 22574 18460 23054
rect 18420 22568 18472 22574
rect 18420 22510 18472 22516
rect 18800 22438 18828 23122
rect 21916 23112 21968 23118
rect 21916 23054 21968 23060
rect 22008 23112 22060 23118
rect 22008 23054 22060 23060
rect 21456 23044 21508 23050
rect 21456 22986 21508 22992
rect 20720 22636 20772 22642
rect 20720 22578 20772 22584
rect 21364 22636 21416 22642
rect 21364 22578 21416 22584
rect 19248 22568 19300 22574
rect 19248 22510 19300 22516
rect 20076 22568 20128 22574
rect 20732 22522 20760 22578
rect 20076 22510 20128 22516
rect 18788 22432 18840 22438
rect 18788 22374 18840 22380
rect 18800 22098 18828 22374
rect 19260 22166 19288 22510
rect 19892 22432 19944 22438
rect 19892 22374 19944 22380
rect 19904 22166 19932 22374
rect 19248 22160 19300 22166
rect 19248 22102 19300 22108
rect 19892 22160 19944 22166
rect 19892 22102 19944 22108
rect 17960 22092 18012 22098
rect 17960 22034 18012 22040
rect 18788 22092 18840 22098
rect 18788 22034 18840 22040
rect 18052 22024 18104 22030
rect 18052 21966 18104 21972
rect 18328 22024 18380 22030
rect 18328 21966 18380 21972
rect 16948 21480 17000 21486
rect 16948 21422 17000 21428
rect 17224 21412 17276 21418
rect 17224 21354 17276 21360
rect 17868 21412 17920 21418
rect 17868 21354 17920 21360
rect 17040 21344 17092 21350
rect 17040 21286 17092 21292
rect 17052 21078 17080 21286
rect 17236 21146 17264 21354
rect 17224 21140 17276 21146
rect 17224 21082 17276 21088
rect 17040 21072 17092 21078
rect 17040 21014 17092 21020
rect 16764 21004 16816 21010
rect 16764 20946 16816 20952
rect 17880 20874 17908 21354
rect 18064 21350 18092 21966
rect 18340 21894 18368 21966
rect 19260 21894 19288 22102
rect 20088 21894 20116 22510
rect 20640 22506 20760 22522
rect 20628 22500 20760 22506
rect 20680 22494 20760 22500
rect 20812 22500 20864 22506
rect 20628 22442 20680 22448
rect 20812 22442 20864 22448
rect 20640 22234 20668 22442
rect 20628 22228 20680 22234
rect 20628 22170 20680 22176
rect 20352 22024 20404 22030
rect 20352 21966 20404 21972
rect 18144 21888 18196 21894
rect 18144 21830 18196 21836
rect 18328 21888 18380 21894
rect 18328 21830 18380 21836
rect 19248 21888 19300 21894
rect 19524 21888 19576 21894
rect 19248 21830 19300 21836
rect 19444 21848 19524 21876
rect 18156 21486 18184 21830
rect 18340 21622 18368 21830
rect 18328 21616 18380 21622
rect 18328 21558 18380 21564
rect 18144 21480 18196 21486
rect 18144 21422 18196 21428
rect 19260 21418 19288 21830
rect 19444 21554 19472 21848
rect 19524 21830 19576 21836
rect 20076 21888 20128 21894
rect 20076 21830 20128 21836
rect 20364 21622 20392 21966
rect 20720 21956 20772 21962
rect 20720 21898 20772 21904
rect 20352 21616 20404 21622
rect 20352 21558 20404 21564
rect 19432 21548 19484 21554
rect 19432 21490 19484 21496
rect 19524 21480 19576 21486
rect 19524 21422 19576 21428
rect 19708 21480 19760 21486
rect 19708 21422 19760 21428
rect 19248 21412 19300 21418
rect 19248 21354 19300 21360
rect 18052 21344 18104 21350
rect 18052 21286 18104 21292
rect 18236 21344 18288 21350
rect 18236 21286 18288 21292
rect 19432 21344 19484 21350
rect 19432 21286 19484 21292
rect 18064 20942 18092 21286
rect 18248 21010 18276 21286
rect 18236 21004 18288 21010
rect 18236 20946 18288 20952
rect 18052 20936 18104 20942
rect 18052 20878 18104 20884
rect 17868 20868 17920 20874
rect 17868 20810 17920 20816
rect 17776 20800 17828 20806
rect 17776 20742 17828 20748
rect 16672 20392 16724 20398
rect 16672 20334 16724 20340
rect 17592 19508 17644 19514
rect 17592 19450 17644 19456
rect 16212 19304 16264 19310
rect 16212 19246 16264 19252
rect 17132 19304 17184 19310
rect 17132 19246 17184 19252
rect 15200 19236 15252 19242
rect 15200 19178 15252 19184
rect 16396 19168 16448 19174
rect 16396 19110 16448 19116
rect 15292 18964 15344 18970
rect 15292 18906 15344 18912
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 14568 18154 14596 18702
rect 15016 18624 15068 18630
rect 15016 18566 15068 18572
rect 14924 18352 14976 18358
rect 14924 18294 14976 18300
rect 14556 18148 14608 18154
rect 14556 18090 14608 18096
rect 14280 17536 14332 17542
rect 14280 17478 14332 17484
rect 14292 17270 14320 17478
rect 14568 17338 14596 18090
rect 14556 17332 14608 17338
rect 14556 17274 14608 17280
rect 14280 17264 14332 17270
rect 14280 17206 14332 17212
rect 14936 15502 14964 18294
rect 15028 18290 15056 18566
rect 15304 18358 15332 18906
rect 15752 18828 15804 18834
rect 15752 18770 15804 18776
rect 15292 18352 15344 18358
rect 15292 18294 15344 18300
rect 15016 18284 15068 18290
rect 15016 18226 15068 18232
rect 15304 18222 15332 18294
rect 15764 18222 15792 18770
rect 16408 18766 16436 19110
rect 17144 18766 17172 19246
rect 17316 19236 17368 19242
rect 17316 19178 17368 19184
rect 17328 18970 17356 19178
rect 17316 18964 17368 18970
rect 17316 18906 17368 18912
rect 17604 18834 17632 19450
rect 17788 19378 17816 20742
rect 19444 20398 19472 21286
rect 19536 21010 19564 21422
rect 19720 21010 19748 21422
rect 20732 21418 20760 21898
rect 20824 21894 20852 22442
rect 21376 22234 21404 22578
rect 21364 22228 21416 22234
rect 21364 22170 21416 22176
rect 21468 22030 21496 22986
rect 21824 22500 21876 22506
rect 21824 22442 21876 22448
rect 21548 22432 21600 22438
rect 21548 22374 21600 22380
rect 21456 22024 21508 22030
rect 21456 21966 21508 21972
rect 20996 21956 21048 21962
rect 20996 21898 21048 21904
rect 21088 21956 21140 21962
rect 21088 21898 21140 21904
rect 20812 21888 20864 21894
rect 20812 21830 20864 21836
rect 20904 21888 20956 21894
rect 20904 21830 20956 21836
rect 20824 21690 20852 21830
rect 20812 21684 20864 21690
rect 20812 21626 20864 21632
rect 20916 21486 20944 21830
rect 21008 21622 21036 21898
rect 20996 21616 21048 21622
rect 20996 21558 21048 21564
rect 21100 21554 21128 21898
rect 21180 21888 21232 21894
rect 21180 21830 21232 21836
rect 21088 21548 21140 21554
rect 21088 21490 21140 21496
rect 20904 21480 20956 21486
rect 20904 21422 20956 21428
rect 20720 21412 20772 21418
rect 20720 21354 20772 21360
rect 20904 21344 20956 21350
rect 21192 21298 21220 21830
rect 21364 21684 21416 21690
rect 21364 21626 21416 21632
rect 21376 21486 21404 21626
rect 21364 21480 21416 21486
rect 21364 21422 21416 21428
rect 20956 21292 21220 21298
rect 20904 21286 21220 21292
rect 20916 21270 21220 21286
rect 19524 21004 19576 21010
rect 19524 20946 19576 20952
rect 19708 21004 19760 21010
rect 19708 20946 19760 20952
rect 20628 21004 20680 21010
rect 20628 20946 20680 20952
rect 19616 20800 19668 20806
rect 19616 20742 19668 20748
rect 19628 20398 19656 20742
rect 20640 20466 20668 20946
rect 20628 20460 20680 20466
rect 20628 20402 20680 20408
rect 19432 20392 19484 20398
rect 19432 20334 19484 20340
rect 19616 20392 19668 20398
rect 19616 20334 19668 20340
rect 20444 20392 20496 20398
rect 20444 20334 20496 20340
rect 19156 20256 19208 20262
rect 19156 20198 19208 20204
rect 19168 19922 19196 20198
rect 18696 19916 18748 19922
rect 18696 19858 18748 19864
rect 19064 19916 19116 19922
rect 19064 19858 19116 19864
rect 19156 19916 19208 19922
rect 19156 19858 19208 19864
rect 19340 19916 19392 19922
rect 19340 19858 19392 19864
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 17788 19242 17816 19314
rect 18708 19310 18736 19858
rect 17960 19304 18012 19310
rect 17960 19246 18012 19252
rect 18696 19304 18748 19310
rect 18696 19246 18748 19252
rect 17776 19236 17828 19242
rect 17776 19178 17828 19184
rect 17788 18902 17816 19178
rect 17972 18970 18000 19246
rect 18420 19236 18472 19242
rect 18420 19178 18472 19184
rect 18052 19168 18104 19174
rect 18052 19110 18104 19116
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 17960 18964 18012 18970
rect 17960 18906 18012 18912
rect 17776 18896 17828 18902
rect 17776 18838 17828 18844
rect 18064 18834 18092 19110
rect 17224 18828 17276 18834
rect 17224 18770 17276 18776
rect 17408 18828 17460 18834
rect 17408 18770 17460 18776
rect 17592 18828 17644 18834
rect 17592 18770 17644 18776
rect 18052 18828 18104 18834
rect 18052 18770 18104 18776
rect 16396 18760 16448 18766
rect 16396 18702 16448 18708
rect 17132 18760 17184 18766
rect 17132 18702 17184 18708
rect 17236 18290 17264 18770
rect 17224 18284 17276 18290
rect 17224 18226 17276 18232
rect 17420 18222 17448 18770
rect 17776 18624 17828 18630
rect 17776 18566 17828 18572
rect 15292 18216 15344 18222
rect 15292 18158 15344 18164
rect 15752 18216 15804 18222
rect 15752 18158 15804 18164
rect 17408 18216 17460 18222
rect 17408 18158 17460 18164
rect 15660 18080 15712 18086
rect 15660 18022 15712 18028
rect 17684 18080 17736 18086
rect 17684 18022 17736 18028
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 15108 16992 15160 16998
rect 15108 16934 15160 16940
rect 15120 16658 15148 16934
rect 15200 16720 15252 16726
rect 15200 16662 15252 16668
rect 15108 16652 15160 16658
rect 15108 16594 15160 16600
rect 15212 15570 15240 16662
rect 15016 15564 15068 15570
rect 15016 15506 15068 15512
rect 15200 15564 15252 15570
rect 15200 15506 15252 15512
rect 14924 15496 14976 15502
rect 14924 15438 14976 15444
rect 14188 14952 14240 14958
rect 14188 14894 14240 14900
rect 15028 14346 15056 15506
rect 15016 14340 15068 14346
rect 15016 14282 15068 14288
rect 14556 13864 14608 13870
rect 14556 13806 14608 13812
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 14292 12986 14320 13126
rect 14280 12980 14332 12986
rect 14280 12922 14332 12928
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 14280 12300 14332 12306
rect 14280 12242 14332 12248
rect 14292 10674 14320 12242
rect 14096 10668 14148 10674
rect 14096 10610 14148 10616
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 13832 9518 13860 10406
rect 13924 9722 13952 10406
rect 14384 10130 14412 12582
rect 14568 12238 14596 13806
rect 14924 12640 14976 12646
rect 14924 12582 14976 12588
rect 14936 12374 14964 12582
rect 14924 12368 14976 12374
rect 14924 12310 14976 12316
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 14924 12096 14976 12102
rect 14924 12038 14976 12044
rect 14936 11762 14964 12038
rect 14924 11756 14976 11762
rect 14924 11698 14976 11704
rect 15028 11626 15056 14282
rect 15304 12850 15332 17818
rect 15672 17202 15700 18022
rect 17696 17746 17724 18022
rect 17788 17746 17816 18566
rect 17684 17740 17736 17746
rect 17684 17682 17736 17688
rect 17776 17740 17828 17746
rect 17776 17682 17828 17688
rect 16764 17264 16816 17270
rect 16764 17206 16816 17212
rect 15660 17196 15712 17202
rect 15660 17138 15712 17144
rect 15384 16788 15436 16794
rect 15384 16730 15436 16736
rect 15396 16046 15424 16730
rect 15672 16658 15700 17138
rect 16028 16992 16080 16998
rect 16028 16934 16080 16940
rect 16040 16726 16068 16934
rect 16028 16720 16080 16726
rect 16028 16662 16080 16668
rect 15660 16652 15712 16658
rect 15660 16594 15712 16600
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15856 16250 15884 16526
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 15936 16244 15988 16250
rect 15936 16186 15988 16192
rect 15948 16130 15976 16186
rect 15672 16102 15976 16130
rect 16040 16114 16068 16662
rect 16488 16448 16540 16454
rect 16488 16390 16540 16396
rect 16028 16108 16080 16114
rect 15384 16040 15436 16046
rect 15384 15982 15436 15988
rect 15396 15570 15424 15982
rect 15384 15564 15436 15570
rect 15384 15506 15436 15512
rect 15672 15366 15700 16102
rect 16028 16050 16080 16056
rect 16500 16046 16528 16390
rect 16776 16046 16804 17206
rect 17788 17202 17816 17682
rect 17868 17536 17920 17542
rect 17868 17478 17920 17484
rect 17776 17196 17828 17202
rect 17776 17138 17828 17144
rect 17880 17134 17908 17478
rect 17868 17128 17920 17134
rect 17868 17070 17920 17076
rect 16856 16788 16908 16794
rect 16856 16730 16908 16736
rect 16868 16250 16896 16730
rect 17880 16658 17908 17070
rect 17960 16992 18012 16998
rect 17960 16934 18012 16940
rect 17132 16652 17184 16658
rect 17132 16594 17184 16600
rect 17316 16652 17368 16658
rect 17316 16594 17368 16600
rect 17868 16652 17920 16658
rect 17868 16594 17920 16600
rect 16948 16584 17000 16590
rect 16948 16526 17000 16532
rect 16856 16244 16908 16250
rect 16856 16186 16908 16192
rect 16960 16046 16988 16526
rect 17144 16046 17172 16594
rect 17328 16250 17356 16594
rect 17972 16250 18000 16934
rect 18156 16794 18184 19110
rect 18432 18970 18460 19178
rect 19076 19174 19104 19858
rect 19168 19310 19196 19858
rect 19156 19304 19208 19310
rect 19156 19246 19208 19252
rect 19064 19168 19116 19174
rect 19064 19110 19116 19116
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 18420 18964 18472 18970
rect 18420 18906 18472 18912
rect 19260 18902 19288 19110
rect 19248 18896 19300 18902
rect 19248 18838 19300 18844
rect 18880 18760 18932 18766
rect 18880 18702 18932 18708
rect 18420 18624 18472 18630
rect 18420 18566 18472 18572
rect 18432 17338 18460 18566
rect 18892 18154 18920 18702
rect 18880 18148 18932 18154
rect 18880 18090 18932 18096
rect 18420 17332 18472 17338
rect 18420 17274 18472 17280
rect 18432 17202 18460 17274
rect 18420 17196 18472 17202
rect 18420 17138 18472 17144
rect 18328 17060 18380 17066
rect 18328 17002 18380 17008
rect 18144 16788 18196 16794
rect 18144 16730 18196 16736
rect 18340 16658 18368 17002
rect 18432 16794 18460 17138
rect 18788 17060 18840 17066
rect 18788 17002 18840 17008
rect 18696 16992 18748 16998
rect 18696 16934 18748 16940
rect 18420 16788 18472 16794
rect 18420 16730 18472 16736
rect 18328 16652 18380 16658
rect 18328 16594 18380 16600
rect 18236 16516 18288 16522
rect 18236 16458 18288 16464
rect 17316 16244 17368 16250
rect 17316 16186 17368 16192
rect 17960 16244 18012 16250
rect 17960 16186 18012 16192
rect 16488 16040 16540 16046
rect 16488 15982 16540 15988
rect 16764 16040 16816 16046
rect 16764 15982 16816 15988
rect 16948 16040 17000 16046
rect 16948 15982 17000 15988
rect 17132 16040 17184 16046
rect 17132 15982 17184 15988
rect 17960 16040 18012 16046
rect 17960 15982 18012 15988
rect 16580 15972 16632 15978
rect 16580 15914 16632 15920
rect 15936 15428 15988 15434
rect 15936 15370 15988 15376
rect 15660 15360 15712 15366
rect 15660 15302 15712 15308
rect 15752 15360 15804 15366
rect 15752 15302 15804 15308
rect 15764 15026 15792 15302
rect 15752 15020 15804 15026
rect 15752 14962 15804 14968
rect 15476 14952 15528 14958
rect 15476 14894 15528 14900
rect 15488 14482 15516 14894
rect 15764 14550 15792 14962
rect 15752 14544 15804 14550
rect 15752 14486 15804 14492
rect 15948 14482 15976 15370
rect 16028 15156 16080 15162
rect 16028 15098 16080 15104
rect 16040 14958 16068 15098
rect 16488 15088 16540 15094
rect 16488 15030 16540 15036
rect 16028 14952 16080 14958
rect 16028 14894 16080 14900
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 16408 14482 16436 14758
rect 16500 14482 16528 15030
rect 16592 14958 16620 15914
rect 16776 14958 16804 15982
rect 17972 15162 18000 15982
rect 18248 15502 18276 16458
rect 18340 15910 18368 16594
rect 18708 16046 18736 16934
rect 18800 16046 18828 17002
rect 18892 16726 18920 18090
rect 18972 17128 19024 17134
rect 18972 17070 19024 17076
rect 19064 17128 19116 17134
rect 19064 17070 19116 17076
rect 18984 16794 19012 17070
rect 18972 16788 19024 16794
rect 18972 16730 19024 16736
rect 18880 16720 18932 16726
rect 18880 16662 18932 16668
rect 18984 16182 19012 16730
rect 18972 16176 19024 16182
rect 18972 16118 19024 16124
rect 18420 16040 18472 16046
rect 18420 15982 18472 15988
rect 18696 16040 18748 16046
rect 18696 15982 18748 15988
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 18328 15904 18380 15910
rect 18328 15846 18380 15852
rect 18236 15496 18288 15502
rect 18236 15438 18288 15444
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 16580 14952 16632 14958
rect 16580 14894 16632 14900
rect 16764 14952 16816 14958
rect 16764 14894 16816 14900
rect 15476 14476 15528 14482
rect 15476 14418 15528 14424
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15936 14476 15988 14482
rect 15936 14418 15988 14424
rect 16396 14476 16448 14482
rect 16396 14418 16448 14424
rect 16488 14476 16540 14482
rect 16488 14418 16540 14424
rect 17776 14476 17828 14482
rect 17776 14418 17828 14424
rect 15384 14272 15436 14278
rect 15384 14214 15436 14220
rect 15396 13870 15424 14214
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15016 11620 15068 11626
rect 15016 11562 15068 11568
rect 15488 11218 15516 14418
rect 15672 14074 15700 14418
rect 17500 14408 17552 14414
rect 17500 14350 17552 14356
rect 16856 14272 16908 14278
rect 16856 14214 16908 14220
rect 15660 14068 15712 14074
rect 15660 14010 15712 14016
rect 16212 14068 16264 14074
rect 16212 14010 16264 14016
rect 15936 12708 15988 12714
rect 15936 12650 15988 12656
rect 15948 12102 15976 12650
rect 15936 12096 15988 12102
rect 15936 12038 15988 12044
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 16132 11694 16160 12038
rect 16224 11898 16252 14010
rect 16868 13870 16896 14214
rect 17512 14074 17540 14350
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 17512 13462 17540 14010
rect 17788 14006 17816 14418
rect 17776 14000 17828 14006
rect 17776 13942 17828 13948
rect 17500 13456 17552 13462
rect 17500 13398 17552 13404
rect 17224 13388 17276 13394
rect 17224 13330 17276 13336
rect 17236 12782 17264 13330
rect 17316 13252 17368 13258
rect 17316 13194 17368 13200
rect 17328 12850 17356 13194
rect 17512 12850 17540 13398
rect 17788 13190 17816 13942
rect 18248 13938 18276 15438
rect 18432 15162 18460 15982
rect 18512 15904 18564 15910
rect 18512 15846 18564 15852
rect 18524 15570 18552 15846
rect 18512 15564 18564 15570
rect 18512 15506 18564 15512
rect 18420 15156 18472 15162
rect 18420 15098 18472 15104
rect 18236 13932 18288 13938
rect 18236 13874 18288 13880
rect 18512 13932 18564 13938
rect 18512 13874 18564 13880
rect 17776 13184 17828 13190
rect 17776 13126 17828 13132
rect 17788 12986 17816 13126
rect 17776 12980 17828 12986
rect 17776 12922 17828 12928
rect 18328 12980 18380 12986
rect 18328 12922 18380 12928
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 17500 12844 17552 12850
rect 17500 12786 17552 12792
rect 17224 12776 17276 12782
rect 17224 12718 17276 12724
rect 16672 12368 16724 12374
rect 16672 12310 16724 12316
rect 16580 12096 16632 12102
rect 16580 12038 16632 12044
rect 16592 11898 16620 12038
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16580 11892 16632 11898
rect 16580 11834 16632 11840
rect 15660 11688 15712 11694
rect 15660 11630 15712 11636
rect 16120 11688 16172 11694
rect 16120 11630 16172 11636
rect 15476 11212 15528 11218
rect 15476 11154 15528 11160
rect 15672 11150 15700 11630
rect 16132 11218 16160 11630
rect 16120 11212 16172 11218
rect 16120 11154 16172 11160
rect 15660 11144 15712 11150
rect 15660 11086 15712 11092
rect 14556 10668 14608 10674
rect 14556 10610 14608 10616
rect 14568 10130 14596 10610
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 14372 10124 14424 10130
rect 14372 10066 14424 10072
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 13912 9716 13964 9722
rect 13912 9658 13964 9664
rect 12900 9512 12952 9518
rect 12900 9454 12952 9460
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 12912 9110 12940 9454
rect 13648 9364 13676 9454
rect 13648 9336 13860 9364
rect 12900 9104 12952 9110
rect 12900 9046 12952 9052
rect 11428 9036 11480 9042
rect 11428 8978 11480 8984
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 10980 8634 11008 8774
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 10980 7954 11008 8570
rect 11152 8560 11204 8566
rect 11152 8502 11204 8508
rect 10968 7948 11020 7954
rect 10968 7890 11020 7896
rect 11164 7886 11192 8502
rect 11440 8430 11468 8978
rect 11612 8968 11664 8974
rect 11612 8910 11664 8916
rect 11624 8430 11652 8910
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12544 8430 12572 8774
rect 12912 8430 12940 9046
rect 13832 8906 13860 9336
rect 13924 8974 13952 9658
rect 13912 8968 13964 8974
rect 13912 8910 13964 8916
rect 14016 8906 14044 10066
rect 15672 9926 15700 11086
rect 15936 11008 15988 11014
rect 15936 10950 15988 10956
rect 15752 10192 15804 10198
rect 15752 10134 15804 10140
rect 14188 9920 14240 9926
rect 14188 9862 14240 9868
rect 15660 9920 15712 9926
rect 15660 9862 15712 9868
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 14108 9042 14136 9318
rect 14096 9036 14148 9042
rect 14096 8978 14148 8984
rect 13820 8900 13872 8906
rect 13820 8842 13872 8848
rect 14004 8900 14056 8906
rect 14004 8842 14056 8848
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 11428 8424 11480 8430
rect 11428 8366 11480 8372
rect 11612 8424 11664 8430
rect 11612 8366 11664 8372
rect 12532 8424 12584 8430
rect 12532 8366 12584 8372
rect 12900 8424 12952 8430
rect 12900 8366 12952 8372
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 11624 7954 11652 8230
rect 11612 7948 11664 7954
rect 11612 7890 11664 7896
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 11612 7744 11664 7750
rect 11612 7686 11664 7692
rect 10692 7336 10744 7342
rect 10692 7278 10744 7284
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 10060 5846 10088 6802
rect 10048 5840 10100 5846
rect 10232 5840 10284 5846
rect 10100 5800 10232 5828
rect 10048 5782 10100 5788
rect 10232 5782 10284 5788
rect 9864 5772 9916 5778
rect 9864 5714 9916 5720
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 8944 5024 8996 5030
rect 8944 4966 8996 4972
rect 8956 4758 8984 4966
rect 8944 4752 8996 4758
rect 8944 4694 8996 4700
rect 8760 4684 8812 4690
rect 8760 4626 8812 4632
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 7196 4480 7248 4486
rect 7196 4422 7248 4428
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 4712 3732 4764 3738
rect 4712 3674 4764 3680
rect 4160 3664 4212 3670
rect 4160 3606 4212 3612
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 3662 3292 3970 3301
rect 3662 3290 3668 3292
rect 3724 3290 3748 3292
rect 3804 3290 3828 3292
rect 3884 3290 3908 3292
rect 3964 3290 3970 3292
rect 3724 3238 3726 3290
rect 3906 3238 3908 3290
rect 3662 3236 3668 3238
rect 3724 3236 3748 3238
rect 3804 3236 3828 3238
rect 3884 3236 3908 3238
rect 3964 3236 3970 3238
rect 3662 3227 3970 3236
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 4172 2990 4200 3606
rect 4816 3602 4844 4014
rect 9416 3942 9444 5102
rect 10060 5030 10088 5782
rect 10704 5778 10732 7278
rect 11072 6798 11100 7686
rect 11624 7410 11652 7686
rect 12820 7410 12848 8230
rect 13556 7954 13584 8434
rect 14108 8430 14136 8978
rect 14200 8838 14228 9862
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 14188 8832 14240 8838
rect 14188 8774 14240 8780
rect 14200 8498 14228 8774
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 14188 8356 14240 8362
rect 14188 8298 14240 8304
rect 14200 8022 14228 8298
rect 15396 8294 15424 9522
rect 15672 9382 15700 9862
rect 15764 9518 15792 10134
rect 15948 10062 15976 10950
rect 16580 10124 16632 10130
rect 16580 10066 16632 10072
rect 15844 10056 15896 10062
rect 15844 9998 15896 10004
rect 15936 10056 15988 10062
rect 15936 9998 15988 10004
rect 15856 9518 15884 9998
rect 16592 9518 16620 10066
rect 16684 9518 16712 12310
rect 17236 12306 17264 12718
rect 17684 12640 17736 12646
rect 17684 12582 17736 12588
rect 17696 12306 17724 12582
rect 17788 12442 17816 12922
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 17960 12708 18012 12714
rect 17960 12650 18012 12656
rect 17776 12436 17828 12442
rect 17776 12378 17828 12384
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 17224 12300 17276 12306
rect 17224 12242 17276 12248
rect 17684 12300 17736 12306
rect 17684 12242 17736 12248
rect 17040 12096 17092 12102
rect 17040 12038 17092 12044
rect 17052 11762 17080 12038
rect 17144 11898 17172 12242
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 17132 11892 17184 11898
rect 17132 11834 17184 11840
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 17328 11694 17356 12038
rect 17316 11688 17368 11694
rect 17316 11630 17368 11636
rect 17972 10266 18000 12650
rect 18064 11898 18092 12786
rect 18144 12776 18196 12782
rect 18144 12718 18196 12724
rect 18236 12776 18288 12782
rect 18236 12718 18288 12724
rect 18156 12374 18184 12718
rect 18248 12442 18276 12718
rect 18340 12442 18368 12922
rect 18236 12436 18288 12442
rect 18236 12378 18288 12384
rect 18328 12436 18380 12442
rect 18328 12378 18380 12384
rect 18144 12368 18196 12374
rect 18144 12310 18196 12316
rect 18052 11892 18104 11898
rect 18052 11834 18104 11840
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 18064 10130 18092 11290
rect 18156 11286 18184 12310
rect 18420 12300 18472 12306
rect 18420 12242 18472 12248
rect 18144 11280 18196 11286
rect 18144 11222 18196 11228
rect 18156 10266 18184 11222
rect 18432 11014 18460 12242
rect 18524 12238 18552 13874
rect 19076 13258 19104 17070
rect 19156 16788 19208 16794
rect 19156 16730 19208 16736
rect 19168 15978 19196 16730
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 19260 16250 19288 16594
rect 19248 16244 19300 16250
rect 19248 16186 19300 16192
rect 19156 15972 19208 15978
rect 19156 15914 19208 15920
rect 19168 14498 19196 15914
rect 19352 14618 19380 19858
rect 19432 19712 19484 19718
rect 19432 19654 19484 19660
rect 19616 19712 19668 19718
rect 19616 19654 19668 19660
rect 20352 19712 20404 19718
rect 20352 19654 20404 19660
rect 19444 19378 19472 19654
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 19628 19310 19656 19654
rect 20364 19446 20392 19654
rect 20352 19440 20404 19446
rect 20352 19382 20404 19388
rect 19616 19304 19668 19310
rect 19616 19246 19668 19252
rect 19708 19304 19760 19310
rect 19708 19246 19760 19252
rect 20352 19304 20404 19310
rect 20352 19246 20404 19252
rect 19628 18834 19656 19246
rect 19616 18828 19668 18834
rect 19616 18770 19668 18776
rect 19628 17202 19656 18770
rect 19720 18426 19748 19246
rect 20364 18970 20392 19246
rect 20456 19242 20484 20334
rect 20640 20330 20668 20402
rect 20720 20392 20772 20398
rect 20772 20340 20852 20346
rect 20720 20334 20852 20340
rect 20628 20324 20680 20330
rect 20732 20318 20852 20334
rect 20628 20266 20680 20272
rect 20720 20256 20772 20262
rect 20720 20198 20772 20204
rect 20536 19712 20588 19718
rect 20536 19654 20588 19660
rect 20548 19310 20576 19654
rect 20536 19304 20588 19310
rect 20536 19246 20588 19252
rect 20444 19236 20496 19242
rect 20444 19178 20496 19184
rect 20352 18964 20404 18970
rect 20352 18906 20404 18912
rect 20076 18624 20128 18630
rect 20076 18566 20128 18572
rect 19708 18420 19760 18426
rect 19708 18362 19760 18368
rect 20088 18222 20116 18566
rect 19892 18216 19944 18222
rect 19892 18158 19944 18164
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 19616 17196 19668 17202
rect 19616 17138 19668 17144
rect 19904 16182 19932 18158
rect 19892 16176 19944 16182
rect 19892 16118 19944 16124
rect 19524 16040 19576 16046
rect 19524 15982 19576 15988
rect 19432 15360 19484 15366
rect 19432 15302 19484 15308
rect 19444 14958 19472 15302
rect 19432 14952 19484 14958
rect 19432 14894 19484 14900
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 19168 14470 19288 14498
rect 19444 14482 19472 14894
rect 19260 14414 19288 14470
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 19248 14408 19300 14414
rect 19248 14350 19300 14356
rect 19444 13938 19472 14418
rect 19432 13932 19484 13938
rect 19432 13874 19484 13880
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 19064 13252 19116 13258
rect 19064 13194 19116 13200
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 18892 12374 18920 12582
rect 18880 12368 18932 12374
rect 18880 12310 18932 12316
rect 18512 12232 18564 12238
rect 18512 12174 18564 12180
rect 19352 11286 19380 13806
rect 19536 12918 19564 15982
rect 20088 14890 20116 18158
rect 20732 17338 20760 20198
rect 20824 19310 20852 20318
rect 20812 19304 20864 19310
rect 20812 19246 20864 19252
rect 20824 18290 20852 19246
rect 20916 18766 20944 21270
rect 20996 20868 21048 20874
rect 20996 20810 21048 20816
rect 21008 20330 21036 20810
rect 21272 20800 21324 20806
rect 21272 20742 21324 20748
rect 20996 20324 21048 20330
rect 20996 20266 21048 20272
rect 21284 20058 21312 20742
rect 21272 20052 21324 20058
rect 21272 19994 21324 20000
rect 20996 19916 21048 19922
rect 20996 19858 21048 19864
rect 20904 18760 20956 18766
rect 20904 18702 20956 18708
rect 21008 18426 21036 19858
rect 21088 19304 21140 19310
rect 21088 19246 21140 19252
rect 21100 18630 21128 19246
rect 21180 19236 21232 19242
rect 21180 19178 21232 19184
rect 21088 18624 21140 18630
rect 21088 18566 21140 18572
rect 20996 18420 21048 18426
rect 20996 18362 21048 18368
rect 20812 18284 20864 18290
rect 20812 18226 20864 18232
rect 20720 17332 20772 17338
rect 20720 17274 20772 17280
rect 20444 17128 20496 17134
rect 20444 17070 20496 17076
rect 20456 16726 20484 17070
rect 20444 16720 20496 16726
rect 20444 16662 20496 16668
rect 21100 15570 21128 18566
rect 21192 18426 21220 19178
rect 21284 18834 21312 19994
rect 21376 19854 21404 21422
rect 21468 21350 21496 21966
rect 21560 21622 21588 22374
rect 21836 22098 21864 22442
rect 21640 22092 21692 22098
rect 21640 22034 21692 22040
rect 21824 22092 21876 22098
rect 21824 22034 21876 22040
rect 21928 22094 21956 23054
rect 22020 22234 22048 23054
rect 22008 22228 22060 22234
rect 22008 22170 22060 22176
rect 22008 22126 22060 22132
rect 21928 22074 22008 22094
rect 21928 22068 22060 22074
rect 22100 22092 22152 22098
rect 21928 22066 22048 22068
rect 21548 21616 21600 21622
rect 21548 21558 21600 21564
rect 21652 21486 21680 22034
rect 21732 21956 21784 21962
rect 21732 21898 21784 21904
rect 21744 21690 21772 21898
rect 21732 21684 21784 21690
rect 21732 21626 21784 21632
rect 21928 21486 21956 22066
rect 22100 22034 22152 22040
rect 22008 22024 22060 22030
rect 22112 21978 22140 22034
rect 22060 21972 22140 21978
rect 22008 21966 22140 21972
rect 22284 22024 22336 22030
rect 22284 21966 22336 21972
rect 22020 21950 22140 21966
rect 22100 21888 22152 21894
rect 22100 21830 22152 21836
rect 21640 21480 21692 21486
rect 21640 21422 21692 21428
rect 21916 21480 21968 21486
rect 21916 21422 21968 21428
rect 21456 21344 21508 21350
rect 21456 21286 21508 21292
rect 21548 20936 21600 20942
rect 21468 20896 21548 20924
rect 21468 20534 21496 20896
rect 21548 20878 21600 20884
rect 21548 20800 21600 20806
rect 21548 20742 21600 20748
rect 21456 20528 21508 20534
rect 21456 20470 21508 20476
rect 21560 20330 21588 20742
rect 21548 20324 21600 20330
rect 21548 20266 21600 20272
rect 21652 19922 21680 21422
rect 21732 21412 21784 21418
rect 21732 21354 21784 21360
rect 21744 21010 21772 21354
rect 21732 21004 21784 21010
rect 21732 20946 21784 20952
rect 22112 20874 22140 21830
rect 22296 21690 22324 21966
rect 22284 21684 22336 21690
rect 22284 21626 22336 21632
rect 22100 20868 22152 20874
rect 22100 20810 22152 20816
rect 21640 19916 21692 19922
rect 21640 19858 21692 19864
rect 21364 19848 21416 19854
rect 21364 19790 21416 19796
rect 21376 19310 21404 19790
rect 23018 19680 23074 19689
rect 23018 19615 23074 19624
rect 23032 19310 23060 19615
rect 21364 19304 21416 19310
rect 21364 19246 21416 19252
rect 21456 19304 21508 19310
rect 21456 19246 21508 19252
rect 22284 19304 22336 19310
rect 22284 19246 22336 19252
rect 22376 19304 22428 19310
rect 22376 19246 22428 19252
rect 22560 19304 22612 19310
rect 22560 19246 22612 19252
rect 23020 19304 23072 19310
rect 23020 19246 23072 19252
rect 21364 19168 21416 19174
rect 21364 19110 21416 19116
rect 21272 18828 21324 18834
rect 21272 18770 21324 18776
rect 21180 18420 21232 18426
rect 21180 18362 21232 18368
rect 21376 18290 21404 19110
rect 21468 18970 21496 19246
rect 21640 19168 21692 19174
rect 21640 19110 21692 19116
rect 21456 18964 21508 18970
rect 21456 18906 21508 18912
rect 21652 18902 21680 19110
rect 21640 18896 21692 18902
rect 21640 18838 21692 18844
rect 22296 18630 22324 19246
rect 21640 18624 21692 18630
rect 21640 18566 21692 18572
rect 22284 18624 22336 18630
rect 22284 18566 22336 18572
rect 21364 18284 21416 18290
rect 21364 18226 21416 18232
rect 21652 18222 21680 18566
rect 22284 18420 22336 18426
rect 22284 18362 22336 18368
rect 21640 18216 21692 18222
rect 21640 18158 21692 18164
rect 22100 17808 22152 17814
rect 22100 17750 22152 17756
rect 21640 17740 21692 17746
rect 21640 17682 21692 17688
rect 22008 17740 22060 17746
rect 22008 17682 22060 17688
rect 21456 16992 21508 16998
rect 21456 16934 21508 16940
rect 21180 16652 21232 16658
rect 21180 16594 21232 16600
rect 21088 15564 21140 15570
rect 21088 15506 21140 15512
rect 20352 15020 20404 15026
rect 20352 14962 20404 14968
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 19892 14884 19944 14890
rect 19892 14826 19944 14832
rect 20076 14884 20128 14890
rect 20076 14826 20128 14832
rect 19904 14482 19932 14826
rect 20364 14482 20392 14962
rect 20628 14884 20680 14890
rect 20628 14826 20680 14832
rect 20640 14482 20668 14826
rect 19892 14476 19944 14482
rect 19892 14418 19944 14424
rect 20352 14476 20404 14482
rect 20352 14418 20404 14424
rect 20628 14476 20680 14482
rect 20628 14418 20680 14424
rect 19616 14272 19668 14278
rect 19616 14214 19668 14220
rect 20168 14272 20220 14278
rect 20168 14214 20220 14220
rect 20812 14272 20864 14278
rect 20812 14214 20864 14220
rect 19628 13938 19656 14214
rect 20180 14074 20208 14214
rect 20168 14068 20220 14074
rect 20168 14010 20220 14016
rect 19616 13932 19668 13938
rect 19616 13874 19668 13880
rect 20824 13870 20852 14214
rect 20916 14074 20944 14962
rect 21088 14612 21140 14618
rect 21088 14554 21140 14560
rect 20904 14068 20956 14074
rect 20904 14010 20956 14016
rect 20812 13864 20864 13870
rect 20812 13806 20864 13812
rect 21100 13802 21128 14554
rect 20168 13796 20220 13802
rect 20168 13738 20220 13744
rect 21088 13796 21140 13802
rect 21088 13738 21140 13744
rect 20180 12986 20208 13738
rect 20720 13728 20772 13734
rect 20720 13670 20772 13676
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 19524 12912 19576 12918
rect 19524 12854 19576 12860
rect 20732 12434 20760 13670
rect 20732 12406 20852 12434
rect 20352 12368 20404 12374
rect 20352 12310 20404 12316
rect 19524 12096 19576 12102
rect 19524 12038 19576 12044
rect 19536 11898 19564 12038
rect 20364 11898 20392 12310
rect 20720 12096 20772 12102
rect 20720 12038 20772 12044
rect 19524 11892 19576 11898
rect 19524 11834 19576 11840
rect 20352 11892 20404 11898
rect 20352 11834 20404 11840
rect 20732 11694 20760 12038
rect 20824 11898 20852 12406
rect 20996 12232 21048 12238
rect 20996 12174 21048 12180
rect 20812 11892 20864 11898
rect 20812 11834 20864 11840
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 19524 11620 19576 11626
rect 19524 11562 19576 11568
rect 19340 11280 19392 11286
rect 19340 11222 19392 11228
rect 19156 11212 19208 11218
rect 19156 11154 19208 11160
rect 19168 11014 19196 11154
rect 19352 11150 19380 11222
rect 19340 11144 19392 11150
rect 19340 11086 19392 11092
rect 18420 11008 18472 11014
rect 18420 10950 18472 10956
rect 19156 11008 19208 11014
rect 19156 10950 19208 10956
rect 18432 10470 18460 10950
rect 18512 10804 18564 10810
rect 18512 10746 18564 10752
rect 18420 10464 18472 10470
rect 18420 10406 18472 10412
rect 18144 10260 18196 10266
rect 18144 10202 18196 10208
rect 16764 10124 16816 10130
rect 16764 10066 16816 10072
rect 18052 10124 18104 10130
rect 18052 10066 18104 10072
rect 15752 9512 15804 9518
rect 15752 9454 15804 9460
rect 15844 9512 15896 9518
rect 15844 9454 15896 9460
rect 16488 9512 16540 9518
rect 16488 9454 16540 9460
rect 16580 9512 16632 9518
rect 16580 9454 16632 9460
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 15660 9376 15712 9382
rect 15660 9318 15712 9324
rect 15672 9178 15700 9318
rect 15660 9172 15712 9178
rect 15660 9114 15712 9120
rect 15568 9036 15620 9042
rect 15568 8978 15620 8984
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 14464 8288 14516 8294
rect 14464 8230 14516 8236
rect 15384 8288 15436 8294
rect 15384 8230 15436 8236
rect 14188 8016 14240 8022
rect 14188 7958 14240 7964
rect 13544 7948 13596 7954
rect 13544 7890 13596 7896
rect 13912 7948 13964 7954
rect 13912 7890 13964 7896
rect 14280 7948 14332 7954
rect 14280 7890 14332 7896
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 13280 7546 13308 7822
rect 13636 7744 13688 7750
rect 13636 7686 13688 7692
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 13648 7410 13676 7686
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 12992 7336 13044 7342
rect 12992 7278 13044 7284
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 11612 7200 11664 7206
rect 11612 7142 11664 7148
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 11164 5914 11192 6802
rect 11624 6662 11652 7142
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 11980 6384 12032 6390
rect 11980 6326 12032 6332
rect 11992 5914 12020 6326
rect 13004 6186 13032 7278
rect 13832 6458 13860 7278
rect 13924 6730 13952 7890
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 14016 7546 14044 7686
rect 14292 7546 14320 7890
rect 14004 7540 14056 7546
rect 14004 7482 14056 7488
rect 14280 7540 14332 7546
rect 14280 7482 14332 7488
rect 14476 7410 14504 8230
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14556 7336 14608 7342
rect 14556 7278 14608 7284
rect 13912 6724 13964 6730
rect 13912 6666 13964 6672
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 14280 6452 14332 6458
rect 14280 6394 14332 6400
rect 12992 6180 13044 6186
rect 12992 6122 13044 6128
rect 13728 6180 13780 6186
rect 13728 6122 13780 6128
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 10692 5772 10744 5778
rect 10692 5714 10744 5720
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 10140 5092 10192 5098
rect 10140 5034 10192 5040
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 10060 4486 10088 4966
rect 10152 4826 10180 5034
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10232 4548 10284 4554
rect 10232 4490 10284 4496
rect 10048 4480 10100 4486
rect 10048 4422 10100 4428
rect 10060 4010 10088 4422
rect 10244 4282 10272 4490
rect 10336 4486 10364 5510
rect 10704 5370 10732 5714
rect 11164 5370 11192 5850
rect 11428 5704 11480 5710
rect 11992 5658 12020 5850
rect 12532 5840 12584 5846
rect 12532 5782 12584 5788
rect 11428 5646 11480 5652
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 10324 4480 10376 4486
rect 10324 4422 10376 4428
rect 10704 4282 10732 5306
rect 10232 4276 10284 4282
rect 10232 4218 10284 4224
rect 10692 4276 10744 4282
rect 10692 4218 10744 4224
rect 10244 4078 10272 4218
rect 11164 4078 11192 5306
rect 11440 5098 11468 5646
rect 11900 5630 12020 5658
rect 11428 5092 11480 5098
rect 11428 5034 11480 5040
rect 11440 4690 11468 5034
rect 11900 4826 11928 5630
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 12072 5568 12124 5574
rect 12072 5510 12124 5516
rect 11888 4820 11940 4826
rect 11888 4762 11940 4768
rect 11428 4684 11480 4690
rect 11428 4626 11480 4632
rect 11992 4146 12020 5510
rect 12084 5166 12112 5510
rect 12072 5160 12124 5166
rect 12072 5102 12124 5108
rect 12544 5098 12572 5782
rect 13004 5778 13032 6122
rect 13360 6112 13412 6118
rect 13360 6054 13412 6060
rect 12992 5772 13044 5778
rect 12992 5714 13044 5720
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 12728 5370 12756 5510
rect 12716 5364 12768 5370
rect 12716 5306 12768 5312
rect 13004 5234 13032 5714
rect 13372 5710 13400 6054
rect 13740 5914 13768 6122
rect 14292 6118 14320 6394
rect 14568 6254 14596 7278
rect 14556 6248 14608 6254
rect 14556 6190 14608 6196
rect 14924 6180 14976 6186
rect 14924 6122 14976 6128
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 14280 6112 14332 6118
rect 14280 6054 14332 6060
rect 14556 6112 14608 6118
rect 14556 6054 14608 6060
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13360 5704 13412 5710
rect 13360 5646 13412 5652
rect 12992 5228 13044 5234
rect 12992 5170 13044 5176
rect 13372 5166 13400 5646
rect 12900 5160 12952 5166
rect 12820 5120 12900 5148
rect 12532 5092 12584 5098
rect 12532 5034 12584 5040
rect 12820 4622 12848 5120
rect 12900 5102 12952 5108
rect 13360 5160 13412 5166
rect 13360 5102 13412 5108
rect 12900 5024 12952 5030
rect 12900 4966 12952 4972
rect 12912 4758 12940 4966
rect 13740 4826 13768 5850
rect 14016 5778 14044 6054
rect 14292 5778 14320 6054
rect 14568 5778 14596 6054
rect 14004 5772 14056 5778
rect 14004 5714 14056 5720
rect 14280 5772 14332 5778
rect 14280 5714 14332 5720
rect 14556 5772 14608 5778
rect 14556 5714 14608 5720
rect 13820 5636 13872 5642
rect 13820 5578 13872 5584
rect 13832 5166 13860 5578
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 14292 5030 14320 5714
rect 14936 5370 14964 6122
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 15212 5574 15240 6054
rect 15396 5846 15424 8230
rect 15488 8090 15516 8570
rect 15580 8362 15608 8978
rect 15752 8900 15804 8906
rect 15752 8842 15804 8848
rect 15764 8430 15792 8842
rect 15752 8424 15804 8430
rect 15752 8366 15804 8372
rect 15568 8356 15620 8362
rect 15568 8298 15620 8304
rect 15476 8084 15528 8090
rect 15476 8026 15528 8032
rect 15568 7336 15620 7342
rect 15568 7278 15620 7284
rect 15580 6934 15608 7278
rect 15764 7154 15792 8366
rect 16212 8356 16264 8362
rect 16212 8298 16264 8304
rect 16224 8090 16252 8298
rect 16212 8084 16264 8090
rect 16212 8026 16264 8032
rect 16500 8022 16528 9454
rect 16592 8650 16620 9454
rect 16684 8906 16712 9454
rect 16672 8900 16724 8906
rect 16672 8842 16724 8848
rect 16592 8634 16712 8650
rect 16592 8628 16724 8634
rect 16592 8622 16672 8628
rect 16672 8570 16724 8576
rect 16488 8016 16540 8022
rect 16488 7958 16540 7964
rect 16500 7342 16528 7958
rect 16684 7886 16712 8570
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 16580 7744 16632 7750
rect 16776 7698 16804 10066
rect 16856 10056 16908 10062
rect 16856 9998 16908 10004
rect 16868 9654 16896 9998
rect 17408 9716 17460 9722
rect 17408 9658 17460 9664
rect 16856 9648 16908 9654
rect 16856 9590 16908 9596
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16868 8090 16896 9318
rect 17420 9178 17448 9658
rect 18064 9518 18092 10066
rect 18156 9586 18184 10202
rect 18432 10130 18460 10406
rect 18524 10266 18552 10746
rect 19168 10742 19196 10950
rect 19352 10810 19380 11086
rect 19536 11014 19564 11562
rect 20824 11506 20852 11834
rect 20732 11478 20852 11506
rect 20628 11280 20680 11286
rect 20628 11222 20680 11228
rect 20640 11150 20668 11222
rect 20732 11150 20760 11478
rect 20628 11144 20680 11150
rect 20628 11086 20680 11092
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 19524 11008 19576 11014
rect 19524 10950 19576 10956
rect 19892 11008 19944 11014
rect 19892 10950 19944 10956
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 19156 10736 19208 10742
rect 19156 10678 19208 10684
rect 19248 10600 19300 10606
rect 19248 10542 19300 10548
rect 18880 10464 18932 10470
rect 18880 10406 18932 10412
rect 18512 10260 18564 10266
rect 18512 10202 18564 10208
rect 18892 10198 18920 10406
rect 18880 10192 18932 10198
rect 18880 10134 18932 10140
rect 18420 10124 18472 10130
rect 18420 10066 18472 10072
rect 18144 9580 18196 9586
rect 18144 9522 18196 9528
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17408 9172 17460 9178
rect 17408 9114 17460 9120
rect 17512 9042 17540 9318
rect 18156 9178 18184 9522
rect 19156 9376 19208 9382
rect 19156 9318 19208 9324
rect 18144 9172 18196 9178
rect 18144 9114 18196 9120
rect 19168 9110 19196 9318
rect 19260 9194 19288 10542
rect 19536 10470 19564 10950
rect 19524 10464 19576 10470
rect 19524 10406 19576 10412
rect 19536 10130 19564 10406
rect 19524 10124 19576 10130
rect 19524 10066 19576 10072
rect 19904 9926 19932 10950
rect 20732 10690 20760 11086
rect 20812 11076 20864 11082
rect 20812 11018 20864 11024
rect 20904 11076 20956 11082
rect 20904 11018 20956 11024
rect 20824 10810 20852 11018
rect 20812 10804 20864 10810
rect 20812 10746 20864 10752
rect 20916 10742 20944 11018
rect 20904 10736 20956 10742
rect 20732 10662 20852 10690
rect 20904 10678 20956 10684
rect 20824 10538 20852 10662
rect 20076 10532 20128 10538
rect 20076 10474 20128 10480
rect 20812 10532 20864 10538
rect 20812 10474 20864 10480
rect 20088 10266 20116 10474
rect 20916 10266 20944 10678
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 20904 10260 20956 10266
rect 20904 10202 20956 10208
rect 20720 10124 20772 10130
rect 20720 10066 20772 10072
rect 19892 9920 19944 9926
rect 19892 9862 19944 9868
rect 20732 9450 20760 10066
rect 20812 9988 20864 9994
rect 20812 9930 20864 9936
rect 20824 9722 20852 9930
rect 20812 9716 20864 9722
rect 20812 9658 20864 9664
rect 20916 9518 20944 10202
rect 21008 10198 21036 12174
rect 21192 11898 21220 16594
rect 21468 16046 21496 16934
rect 21652 16250 21680 17682
rect 21732 17536 21784 17542
rect 21732 17478 21784 17484
rect 21744 16658 21772 17478
rect 21732 16652 21784 16658
rect 21732 16594 21784 16600
rect 22020 16250 22048 17682
rect 21640 16244 21692 16250
rect 21640 16186 21692 16192
rect 22008 16244 22060 16250
rect 22008 16186 22060 16192
rect 21456 16040 21508 16046
rect 21456 15982 21508 15988
rect 21548 16040 21600 16046
rect 21548 15982 21600 15988
rect 21468 15434 21496 15982
rect 21560 15638 21588 15982
rect 21732 15904 21784 15910
rect 21732 15846 21784 15852
rect 21548 15632 21600 15638
rect 21548 15574 21600 15580
rect 21456 15428 21508 15434
rect 21376 15388 21456 15416
rect 21376 14958 21404 15388
rect 21456 15370 21508 15376
rect 21560 15162 21588 15574
rect 21548 15156 21600 15162
rect 21548 15098 21600 15104
rect 21456 15020 21508 15026
rect 21456 14962 21508 14968
rect 21364 14952 21416 14958
rect 21364 14894 21416 14900
rect 21468 13938 21496 14962
rect 21456 13932 21508 13938
rect 21456 13874 21508 13880
rect 21548 13864 21600 13870
rect 21548 13806 21600 13812
rect 21456 13388 21508 13394
rect 21456 13330 21508 13336
rect 21180 11892 21232 11898
rect 21180 11834 21232 11840
rect 21180 10600 21232 10606
rect 21180 10542 21232 10548
rect 20996 10192 21048 10198
rect 20996 10134 21048 10140
rect 20904 9512 20956 9518
rect 20904 9454 20956 9460
rect 20720 9444 20772 9450
rect 20720 9386 20772 9392
rect 19260 9178 19380 9194
rect 19260 9172 19392 9178
rect 19260 9166 19340 9172
rect 19156 9104 19208 9110
rect 19156 9046 19208 9052
rect 17500 9036 17552 9042
rect 17500 8978 17552 8984
rect 19156 8288 19208 8294
rect 19156 8230 19208 8236
rect 16856 8084 16908 8090
rect 16856 8026 16908 8032
rect 16868 7954 16896 8026
rect 16856 7948 16908 7954
rect 16856 7890 16908 7896
rect 18328 7948 18380 7954
rect 18328 7890 18380 7896
rect 18788 7948 18840 7954
rect 18788 7890 18840 7896
rect 16632 7692 16804 7698
rect 16580 7686 16804 7692
rect 16592 7670 16804 7686
rect 16868 7410 16896 7890
rect 16856 7404 16908 7410
rect 16856 7346 16908 7352
rect 16488 7336 16540 7342
rect 16488 7278 16540 7284
rect 16212 7200 16264 7206
rect 15764 7126 15976 7154
rect 16212 7142 16264 7148
rect 15568 6928 15620 6934
rect 15568 6870 15620 6876
rect 15580 6458 15608 6870
rect 15948 6798 15976 7126
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 15568 6452 15620 6458
rect 15568 6394 15620 6400
rect 15384 5840 15436 5846
rect 15384 5782 15436 5788
rect 15580 5778 15608 6394
rect 15948 6118 15976 6734
rect 16120 6656 16172 6662
rect 16120 6598 16172 6604
rect 16132 6186 16160 6598
rect 16224 6458 16252 7142
rect 16500 6934 16528 7278
rect 16488 6928 16540 6934
rect 16488 6870 16540 6876
rect 18340 6866 18368 7890
rect 18800 7546 18828 7890
rect 18788 7540 18840 7546
rect 18788 7482 18840 7488
rect 19168 7274 19196 8230
rect 19260 8022 19288 9166
rect 19340 9114 19392 9120
rect 20812 8968 20864 8974
rect 20812 8910 20864 8916
rect 20824 8838 20852 8910
rect 20812 8832 20864 8838
rect 20812 8774 20864 8780
rect 19248 8016 19300 8022
rect 19248 7958 19300 7964
rect 19892 7812 19944 7818
rect 19892 7754 19944 7760
rect 19904 7410 19932 7754
rect 20720 7540 20772 7546
rect 20720 7482 20772 7488
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 19892 7404 19944 7410
rect 19892 7346 19944 7352
rect 19156 7268 19208 7274
rect 19156 7210 19208 7216
rect 16396 6860 16448 6866
rect 16396 6802 16448 6808
rect 18328 6860 18380 6866
rect 18328 6802 18380 6808
rect 18604 6860 18656 6866
rect 18604 6802 18656 6808
rect 16408 6458 16436 6802
rect 16212 6452 16264 6458
rect 16212 6394 16264 6400
rect 16396 6452 16448 6458
rect 16396 6394 16448 6400
rect 16028 6180 16080 6186
rect 16028 6122 16080 6128
rect 16120 6180 16172 6186
rect 16120 6122 16172 6128
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 16040 5846 16068 6122
rect 16488 6112 16540 6118
rect 16488 6054 16540 6060
rect 16028 5840 16080 5846
rect 16028 5782 16080 5788
rect 15568 5772 15620 5778
rect 15568 5714 15620 5720
rect 15200 5568 15252 5574
rect 15200 5510 15252 5516
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 14924 5364 14976 5370
rect 14924 5306 14976 5312
rect 15396 5166 15424 5510
rect 16500 5234 16528 6054
rect 18340 5778 18368 6802
rect 18616 6458 18644 6802
rect 19168 6458 19196 7210
rect 19340 7200 19392 7206
rect 19340 7142 19392 7148
rect 18604 6452 18656 6458
rect 18604 6394 18656 6400
rect 19156 6452 19208 6458
rect 19156 6394 19208 6400
rect 18328 5772 18380 5778
rect 18328 5714 18380 5720
rect 18880 5772 18932 5778
rect 18880 5714 18932 5720
rect 18892 5370 18920 5714
rect 19168 5370 19196 6394
rect 19352 6254 19380 7142
rect 19444 6458 19472 7346
rect 19800 7336 19852 7342
rect 19800 7278 19852 7284
rect 19708 6724 19760 6730
rect 19708 6666 19760 6672
rect 19432 6452 19484 6458
rect 19432 6394 19484 6400
rect 19444 6322 19472 6394
rect 19720 6322 19748 6666
rect 19812 6458 19840 7278
rect 19904 6866 19932 7346
rect 19984 7268 20036 7274
rect 19984 7210 20036 7216
rect 19996 6934 20024 7210
rect 20536 7200 20588 7206
rect 20536 7142 20588 7148
rect 19984 6928 20036 6934
rect 19984 6870 20036 6876
rect 19892 6860 19944 6866
rect 19892 6802 19944 6808
rect 20260 6860 20312 6866
rect 20260 6802 20312 6808
rect 19984 6656 20036 6662
rect 19984 6598 20036 6604
rect 19996 6458 20024 6598
rect 19800 6452 19852 6458
rect 19800 6394 19852 6400
rect 19984 6452 20036 6458
rect 19984 6394 20036 6400
rect 19432 6316 19484 6322
rect 19432 6258 19484 6264
rect 19708 6316 19760 6322
rect 19708 6258 19760 6264
rect 19812 6254 19840 6394
rect 19340 6248 19392 6254
rect 19340 6190 19392 6196
rect 19800 6248 19852 6254
rect 19800 6190 19852 6196
rect 19708 5840 19760 5846
rect 19708 5782 19760 5788
rect 18880 5364 18932 5370
rect 18880 5306 18932 5312
rect 19156 5364 19208 5370
rect 19156 5306 19208 5312
rect 16488 5228 16540 5234
rect 16488 5170 16540 5176
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 14280 5024 14332 5030
rect 14280 4966 14332 4972
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 12900 4752 12952 4758
rect 12900 4694 12952 4700
rect 19720 4622 19748 5782
rect 19812 5302 19840 6190
rect 19996 5914 20024 6394
rect 20272 6186 20300 6802
rect 20548 6322 20576 7142
rect 20732 6730 20760 7482
rect 20720 6724 20772 6730
rect 20720 6666 20772 6672
rect 20536 6316 20588 6322
rect 20536 6258 20588 6264
rect 20260 6180 20312 6186
rect 20260 6122 20312 6128
rect 20272 5914 20300 6122
rect 20548 6066 20576 6258
rect 20548 6038 20668 6066
rect 19984 5908 20036 5914
rect 19984 5850 20036 5856
rect 20260 5908 20312 5914
rect 20260 5850 20312 5856
rect 20076 5568 20128 5574
rect 20076 5510 20128 5516
rect 19800 5296 19852 5302
rect 19800 5238 19852 5244
rect 20088 5098 20116 5510
rect 20272 5166 20300 5850
rect 20640 5778 20668 6038
rect 20352 5772 20404 5778
rect 20352 5714 20404 5720
rect 20628 5772 20680 5778
rect 20628 5714 20680 5720
rect 20364 5166 20392 5714
rect 20260 5160 20312 5166
rect 20260 5102 20312 5108
rect 20352 5160 20404 5166
rect 20640 5148 20668 5714
rect 20732 5710 20760 6666
rect 20824 6186 20852 8774
rect 21008 8362 21036 10134
rect 21192 9586 21220 10542
rect 21272 9920 21324 9926
rect 21272 9862 21324 9868
rect 21364 9920 21416 9926
rect 21364 9862 21416 9868
rect 21180 9580 21232 9586
rect 21180 9522 21232 9528
rect 20996 8356 21048 8362
rect 20996 8298 21048 8304
rect 20996 7336 21048 7342
rect 20996 7278 21048 7284
rect 20904 6792 20956 6798
rect 20904 6734 20956 6740
rect 20916 6458 20944 6734
rect 20904 6452 20956 6458
rect 20904 6394 20956 6400
rect 20812 6180 20864 6186
rect 20812 6122 20864 6128
rect 20720 5704 20772 5710
rect 20720 5646 20772 5652
rect 20824 5370 20852 6122
rect 21008 5914 21036 7278
rect 21192 6866 21220 9522
rect 21284 9450 21312 9862
rect 21376 9722 21404 9862
rect 21364 9716 21416 9722
rect 21364 9658 21416 9664
rect 21272 9444 21324 9450
rect 21272 9386 21324 9392
rect 21364 9036 21416 9042
rect 21364 8978 21416 8984
rect 21376 8634 21404 8978
rect 21364 8628 21416 8634
rect 21364 8570 21416 8576
rect 21272 8356 21324 8362
rect 21272 8298 21324 8304
rect 21284 7206 21312 8298
rect 21468 8090 21496 13330
rect 21560 12434 21588 13806
rect 21744 13462 21772 15846
rect 22020 15722 22048 16186
rect 22112 16046 22140 17750
rect 22192 17060 22244 17066
rect 22192 17002 22244 17008
rect 22204 16114 22232 17002
rect 22296 16182 22324 18362
rect 22388 17134 22416 19246
rect 22376 17128 22428 17134
rect 22376 17070 22428 17076
rect 22284 16176 22336 16182
rect 22284 16118 22336 16124
rect 22192 16108 22244 16114
rect 22192 16050 22244 16056
rect 22100 16040 22152 16046
rect 22100 15982 22152 15988
rect 21824 15700 21876 15706
rect 21824 15642 21876 15648
rect 21928 15694 22048 15722
rect 21836 15502 21864 15642
rect 21824 15496 21876 15502
rect 21824 15438 21876 15444
rect 21836 14890 21864 15438
rect 21824 14884 21876 14890
rect 21824 14826 21876 14832
rect 21732 13456 21784 13462
rect 21652 13416 21732 13444
rect 21652 12918 21680 13416
rect 21732 13398 21784 13404
rect 21732 13320 21784 13326
rect 21732 13262 21784 13268
rect 21744 12986 21772 13262
rect 21732 12980 21784 12986
rect 21732 12922 21784 12928
rect 21640 12912 21692 12918
rect 21640 12854 21692 12860
rect 21836 12850 21864 14826
rect 21928 13530 21956 15694
rect 22008 15564 22060 15570
rect 22008 15506 22060 15512
rect 22020 14958 22048 15506
rect 22296 15366 22324 16118
rect 22468 15428 22520 15434
rect 22468 15370 22520 15376
rect 22284 15360 22336 15366
rect 22284 15302 22336 15308
rect 22008 14952 22060 14958
rect 22008 14894 22060 14900
rect 22008 14068 22060 14074
rect 22008 14010 22060 14016
rect 21916 13524 21968 13530
rect 21916 13466 21968 13472
rect 21824 12844 21876 12850
rect 21824 12786 21876 12792
rect 21560 12406 21680 12434
rect 21548 12300 21600 12306
rect 21548 12242 21600 12248
rect 21560 12170 21588 12242
rect 21548 12164 21600 12170
rect 21548 12106 21600 12112
rect 21560 11286 21588 12106
rect 21652 11898 21680 12406
rect 21928 12306 21956 13466
rect 22020 13190 22048 14010
rect 22480 13870 22508 15370
rect 22572 14890 22600 19246
rect 22652 18760 22704 18766
rect 22652 18702 22704 18708
rect 22664 16726 22692 18702
rect 22836 17808 22888 17814
rect 22836 17750 22888 17756
rect 22848 17338 22876 17750
rect 22836 17332 22888 17338
rect 22836 17274 22888 17280
rect 22836 17128 22888 17134
rect 22836 17070 22888 17076
rect 22744 16992 22796 16998
rect 22744 16934 22796 16940
rect 22652 16720 22704 16726
rect 22652 16662 22704 16668
rect 22560 14884 22612 14890
rect 22560 14826 22612 14832
rect 22468 13864 22520 13870
rect 22468 13806 22520 13812
rect 22560 13796 22612 13802
rect 22560 13738 22612 13744
rect 22284 13456 22336 13462
rect 22284 13398 22336 13404
rect 22192 13252 22244 13258
rect 22192 13194 22244 13200
rect 22008 13184 22060 13190
rect 22008 13126 22060 13132
rect 22204 12646 22232 13194
rect 22192 12640 22244 12646
rect 22192 12582 22244 12588
rect 21916 12300 21968 12306
rect 21916 12242 21968 12248
rect 22100 12300 22152 12306
rect 22100 12242 22152 12248
rect 22008 12096 22060 12102
rect 22008 12038 22060 12044
rect 21640 11892 21692 11898
rect 21640 11834 21692 11840
rect 21548 11280 21600 11286
rect 21548 11222 21600 11228
rect 21560 10198 21588 11222
rect 21652 10810 21680 11834
rect 21824 11620 21876 11626
rect 21824 11562 21876 11568
rect 21836 11354 21864 11562
rect 21824 11348 21876 11354
rect 21824 11290 21876 11296
rect 22020 11286 22048 12038
rect 22008 11280 22060 11286
rect 22008 11222 22060 11228
rect 22112 11082 22140 12242
rect 22100 11076 22152 11082
rect 22100 11018 22152 11024
rect 21640 10804 21692 10810
rect 21640 10746 21692 10752
rect 21548 10192 21600 10198
rect 21548 10134 21600 10140
rect 22008 9988 22060 9994
rect 22008 9930 22060 9936
rect 21916 9920 21968 9926
rect 21916 9862 21968 9868
rect 21928 8566 21956 9862
rect 22020 8634 22048 9930
rect 22008 8628 22060 8634
rect 22008 8570 22060 8576
rect 21916 8560 21968 8566
rect 21916 8502 21968 8508
rect 21456 8084 21508 8090
rect 21456 8026 21508 8032
rect 21824 8016 21876 8022
rect 21824 7958 21876 7964
rect 21456 7880 21508 7886
rect 21456 7822 21508 7828
rect 21364 7744 21416 7750
rect 21364 7686 21416 7692
rect 21376 7546 21404 7686
rect 21364 7540 21416 7546
rect 21364 7482 21416 7488
rect 21272 7200 21324 7206
rect 21272 7142 21324 7148
rect 21180 6860 21232 6866
rect 21180 6802 21232 6808
rect 21192 6338 21220 6802
rect 21284 6798 21312 7142
rect 21468 7002 21496 7822
rect 21836 7274 21864 7958
rect 21928 7954 21956 8502
rect 21916 7948 21968 7954
rect 21916 7890 21968 7896
rect 21928 7410 21956 7890
rect 21916 7404 21968 7410
rect 21916 7346 21968 7352
rect 21824 7268 21876 7274
rect 21824 7210 21876 7216
rect 21548 7200 21600 7206
rect 21548 7142 21600 7148
rect 21456 6996 21508 7002
rect 21456 6938 21508 6944
rect 21560 6934 21588 7142
rect 21548 6928 21600 6934
rect 21548 6870 21600 6876
rect 21272 6792 21324 6798
rect 21272 6734 21324 6740
rect 21836 6662 21864 7210
rect 21272 6656 21324 6662
rect 21272 6598 21324 6604
rect 21824 6656 21876 6662
rect 21824 6598 21876 6604
rect 21100 6310 21220 6338
rect 21100 6254 21128 6310
rect 21088 6248 21140 6254
rect 21088 6190 21140 6196
rect 20996 5908 21048 5914
rect 20996 5850 21048 5856
rect 21284 5778 21312 6598
rect 21836 5778 21864 6598
rect 21928 5778 21956 7346
rect 22112 6458 22140 11018
rect 22204 10198 22232 12582
rect 22192 10192 22244 10198
rect 22192 10134 22244 10140
rect 22192 7404 22244 7410
rect 22192 7346 22244 7352
rect 22100 6452 22152 6458
rect 22100 6394 22152 6400
rect 21272 5772 21324 5778
rect 21272 5714 21324 5720
rect 21824 5772 21876 5778
rect 21824 5714 21876 5720
rect 21916 5772 21968 5778
rect 21916 5714 21968 5720
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 22204 5166 22232 7346
rect 22296 5642 22324 13398
rect 22468 13388 22520 13394
rect 22468 13330 22520 13336
rect 22480 12714 22508 13330
rect 22468 12708 22520 12714
rect 22468 12650 22520 12656
rect 22376 11688 22428 11694
rect 22376 11630 22428 11636
rect 22388 7410 22416 11630
rect 22572 10198 22600 13738
rect 22756 12442 22784 16934
rect 22848 16794 22876 17070
rect 22836 16788 22888 16794
rect 22836 16730 22888 16736
rect 22836 14884 22888 14890
rect 22836 14826 22888 14832
rect 22848 13326 22876 14826
rect 22836 13320 22888 13326
rect 22836 13262 22888 13268
rect 22744 12436 22796 12442
rect 22744 12378 22796 12384
rect 22468 10192 22520 10198
rect 22468 10134 22520 10140
rect 22560 10192 22612 10198
rect 22560 10134 22612 10140
rect 22480 9722 22508 10134
rect 22572 9926 22600 10134
rect 22560 9920 22612 9926
rect 22560 9862 22612 9868
rect 22468 9716 22520 9722
rect 22468 9658 22520 9664
rect 22480 9382 22508 9658
rect 22468 9376 22520 9382
rect 22468 9318 22520 9324
rect 22572 9178 22600 9862
rect 22560 9172 22612 9178
rect 22560 9114 22612 9120
rect 22848 7886 22876 13262
rect 23020 12300 23072 12306
rect 23020 12242 23072 12248
rect 23032 11801 23060 12242
rect 23018 11792 23074 11801
rect 23018 11727 23074 11736
rect 22836 7880 22888 7886
rect 22836 7822 22888 7828
rect 22376 7404 22428 7410
rect 22376 7346 22428 7352
rect 22468 7336 22520 7342
rect 22468 7278 22520 7284
rect 22284 5636 22336 5642
rect 22284 5578 22336 5584
rect 20720 5160 20772 5166
rect 20640 5120 20720 5148
rect 20352 5102 20404 5108
rect 20720 5102 20772 5108
rect 20904 5160 20956 5166
rect 20904 5102 20956 5108
rect 22192 5160 22244 5166
rect 22192 5102 22244 5108
rect 20076 5092 20128 5098
rect 20076 5034 20128 5040
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 19996 4758 20024 4966
rect 20272 4826 20300 5102
rect 20916 4826 20944 5102
rect 20260 4820 20312 4826
rect 20260 4762 20312 4768
rect 20904 4820 20956 4826
rect 20904 4762 20956 4768
rect 19984 4752 20036 4758
rect 19984 4694 20036 4700
rect 12808 4616 12860 4622
rect 12808 4558 12860 4564
rect 19708 4616 19760 4622
rect 19708 4558 19760 4564
rect 22480 4486 22508 7278
rect 22560 6248 22612 6254
rect 22560 6190 22612 6196
rect 22572 5914 22600 6190
rect 22836 6112 22888 6118
rect 22836 6054 22888 6060
rect 22560 5908 22612 5914
rect 22560 5850 22612 5856
rect 22848 5778 22876 6054
rect 22836 5772 22888 5778
rect 22836 5714 22888 5720
rect 22468 4480 22520 4486
rect 22468 4422 22520 4428
rect 22836 4480 22888 4486
rect 22836 4422 22888 4428
rect 22848 4282 22876 4422
rect 22836 4276 22888 4282
rect 22836 4218 22888 4224
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 10232 4072 10284 4078
rect 10232 4014 10284 4020
rect 11152 4072 11204 4078
rect 11152 4014 11204 4020
rect 23020 4072 23072 4078
rect 23020 4014 23072 4020
rect 10048 4004 10100 4010
rect 10048 3946 10100 3952
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 9404 3936 9456 3942
rect 23032 3913 23060 4014
rect 9404 3878 9456 3884
rect 23018 3904 23074 3913
rect 5460 3670 5488 3878
rect 23018 3839 23074 3848
rect 5448 3664 5500 3670
rect 5448 3606 5500 3612
rect 4804 3596 4856 3602
rect 4804 3538 4856 3544
rect 3148 2984 3200 2990
rect 3148 2926 3200 2932
rect 4160 2984 4212 2990
rect 4160 2926 4212 2932
rect 4322 2748 4630 2757
rect 4322 2746 4328 2748
rect 4384 2746 4408 2748
rect 4464 2746 4488 2748
rect 4544 2746 4568 2748
rect 4624 2746 4630 2748
rect 4384 2694 4386 2746
rect 4566 2694 4568 2746
rect 4322 2692 4328 2694
rect 4384 2692 4408 2694
rect 4464 2692 4488 2694
rect 4544 2692 4568 2694
rect 4624 2692 4630 2694
rect 4322 2683 4630 2692
rect 3662 2204 3970 2213
rect 3662 2202 3668 2204
rect 3724 2202 3748 2204
rect 3804 2202 3828 2204
rect 3884 2202 3908 2204
rect 3964 2202 3970 2204
rect 3724 2150 3726 2202
rect 3906 2150 3908 2202
rect 3662 2148 3668 2150
rect 3724 2148 3748 2150
rect 3804 2148 3828 2150
rect 3884 2148 3908 2150
rect 3964 2148 3970 2150
rect 3662 2139 3970 2148
rect 4322 1660 4630 1669
rect 4322 1658 4328 1660
rect 4384 1658 4408 1660
rect 4464 1658 4488 1660
rect 4544 1658 4568 1660
rect 4624 1658 4630 1660
rect 4384 1606 4386 1658
rect 4566 1606 4568 1658
rect 4322 1604 4328 1606
rect 4384 1604 4408 1606
rect 4464 1604 4488 1606
rect 4544 1604 4568 1606
rect 4624 1604 4630 1606
rect 4322 1595 4630 1604
rect 3662 1116 3970 1125
rect 3662 1114 3668 1116
rect 3724 1114 3748 1116
rect 3804 1114 3828 1116
rect 3884 1114 3908 1116
rect 3964 1114 3970 1116
rect 3724 1062 3726 1114
rect 3906 1062 3908 1114
rect 3662 1060 3668 1062
rect 3724 1060 3748 1062
rect 3804 1060 3828 1062
rect 3884 1060 3908 1062
rect 3964 1060 3970 1062
rect 3662 1051 3970 1060
rect 4322 572 4630 581
rect 4322 570 4328 572
rect 4384 570 4408 572
rect 4464 570 4488 572
rect 4544 570 4568 572
rect 4624 570 4630 572
rect 4384 518 4386 570
rect 4566 518 4568 570
rect 4322 516 4328 518
rect 4384 516 4408 518
rect 4464 516 4488 518
rect 4544 516 4568 518
rect 4624 516 4630 518
rect 4322 507 4630 516
<< via2 >>
rect 4328 23418 4384 23420
rect 4408 23418 4464 23420
rect 4488 23418 4544 23420
rect 4568 23418 4624 23420
rect 4328 23366 4374 23418
rect 4374 23366 4384 23418
rect 4408 23366 4438 23418
rect 4438 23366 4450 23418
rect 4450 23366 4464 23418
rect 4488 23366 4502 23418
rect 4502 23366 4514 23418
rect 4514 23366 4544 23418
rect 4568 23366 4578 23418
rect 4578 23366 4624 23418
rect 4328 23364 4384 23366
rect 4408 23364 4464 23366
rect 4488 23364 4544 23366
rect 4568 23364 4624 23366
rect 3668 22874 3724 22876
rect 3748 22874 3804 22876
rect 3828 22874 3884 22876
rect 3908 22874 3964 22876
rect 3668 22822 3714 22874
rect 3714 22822 3724 22874
rect 3748 22822 3778 22874
rect 3778 22822 3790 22874
rect 3790 22822 3804 22874
rect 3828 22822 3842 22874
rect 3842 22822 3854 22874
rect 3854 22822 3884 22874
rect 3908 22822 3918 22874
rect 3918 22822 3964 22874
rect 3668 22820 3724 22822
rect 3748 22820 3804 22822
rect 3828 22820 3884 22822
rect 3908 22820 3964 22822
rect 4328 22330 4384 22332
rect 4408 22330 4464 22332
rect 4488 22330 4544 22332
rect 4568 22330 4624 22332
rect 4328 22278 4374 22330
rect 4374 22278 4384 22330
rect 4408 22278 4438 22330
rect 4438 22278 4450 22330
rect 4450 22278 4464 22330
rect 4488 22278 4502 22330
rect 4502 22278 4514 22330
rect 4514 22278 4544 22330
rect 4568 22278 4578 22330
rect 4578 22278 4624 22330
rect 4328 22276 4384 22278
rect 4408 22276 4464 22278
rect 4488 22276 4544 22278
rect 4568 22276 4624 22278
rect 3668 21786 3724 21788
rect 3748 21786 3804 21788
rect 3828 21786 3884 21788
rect 3908 21786 3964 21788
rect 3668 21734 3714 21786
rect 3714 21734 3724 21786
rect 3748 21734 3778 21786
rect 3778 21734 3790 21786
rect 3790 21734 3804 21786
rect 3828 21734 3842 21786
rect 3842 21734 3854 21786
rect 3854 21734 3884 21786
rect 3908 21734 3918 21786
rect 3918 21734 3964 21786
rect 3668 21732 3724 21734
rect 3748 21732 3804 21734
rect 3828 21732 3884 21734
rect 3908 21732 3964 21734
rect 4328 21242 4384 21244
rect 4408 21242 4464 21244
rect 4488 21242 4544 21244
rect 4568 21242 4624 21244
rect 4328 21190 4374 21242
rect 4374 21190 4384 21242
rect 4408 21190 4438 21242
rect 4438 21190 4450 21242
rect 4450 21190 4464 21242
rect 4488 21190 4502 21242
rect 4502 21190 4514 21242
rect 4514 21190 4544 21242
rect 4568 21190 4578 21242
rect 4578 21190 4624 21242
rect 4328 21188 4384 21190
rect 4408 21188 4464 21190
rect 4488 21188 4544 21190
rect 4568 21188 4624 21190
rect 3668 20698 3724 20700
rect 3748 20698 3804 20700
rect 3828 20698 3884 20700
rect 3908 20698 3964 20700
rect 3668 20646 3714 20698
rect 3714 20646 3724 20698
rect 3748 20646 3778 20698
rect 3778 20646 3790 20698
rect 3790 20646 3804 20698
rect 3828 20646 3842 20698
rect 3842 20646 3854 20698
rect 3854 20646 3884 20698
rect 3908 20646 3918 20698
rect 3918 20646 3964 20698
rect 3668 20644 3724 20646
rect 3748 20644 3804 20646
rect 3828 20644 3884 20646
rect 3908 20644 3964 20646
rect 4328 20154 4384 20156
rect 4408 20154 4464 20156
rect 4488 20154 4544 20156
rect 4568 20154 4624 20156
rect 4328 20102 4374 20154
rect 4374 20102 4384 20154
rect 4408 20102 4438 20154
rect 4438 20102 4450 20154
rect 4450 20102 4464 20154
rect 4488 20102 4502 20154
rect 4502 20102 4514 20154
rect 4514 20102 4544 20154
rect 4568 20102 4578 20154
rect 4578 20102 4624 20154
rect 4328 20100 4384 20102
rect 4408 20100 4464 20102
rect 4488 20100 4544 20102
rect 4568 20100 4624 20102
rect 3668 19610 3724 19612
rect 3748 19610 3804 19612
rect 3828 19610 3884 19612
rect 3908 19610 3964 19612
rect 3668 19558 3714 19610
rect 3714 19558 3724 19610
rect 3748 19558 3778 19610
rect 3778 19558 3790 19610
rect 3790 19558 3804 19610
rect 3828 19558 3842 19610
rect 3842 19558 3854 19610
rect 3854 19558 3884 19610
rect 3908 19558 3918 19610
rect 3918 19558 3964 19610
rect 3668 19556 3724 19558
rect 3748 19556 3804 19558
rect 3828 19556 3884 19558
rect 3908 19556 3964 19558
rect 3668 18522 3724 18524
rect 3748 18522 3804 18524
rect 3828 18522 3884 18524
rect 3908 18522 3964 18524
rect 3668 18470 3714 18522
rect 3714 18470 3724 18522
rect 3748 18470 3778 18522
rect 3778 18470 3790 18522
rect 3790 18470 3804 18522
rect 3828 18470 3842 18522
rect 3842 18470 3854 18522
rect 3854 18470 3884 18522
rect 3908 18470 3918 18522
rect 3918 18470 3964 18522
rect 3668 18468 3724 18470
rect 3748 18468 3804 18470
rect 3828 18468 3884 18470
rect 3908 18468 3964 18470
rect 3668 17434 3724 17436
rect 3748 17434 3804 17436
rect 3828 17434 3884 17436
rect 3908 17434 3964 17436
rect 3668 17382 3714 17434
rect 3714 17382 3724 17434
rect 3748 17382 3778 17434
rect 3778 17382 3790 17434
rect 3790 17382 3804 17434
rect 3828 17382 3842 17434
rect 3842 17382 3854 17434
rect 3854 17382 3884 17434
rect 3908 17382 3918 17434
rect 3918 17382 3964 17434
rect 3668 17380 3724 17382
rect 3748 17380 3804 17382
rect 3828 17380 3884 17382
rect 3908 17380 3964 17382
rect 4328 19066 4384 19068
rect 4408 19066 4464 19068
rect 4488 19066 4544 19068
rect 4568 19066 4624 19068
rect 4328 19014 4374 19066
rect 4374 19014 4384 19066
rect 4408 19014 4438 19066
rect 4438 19014 4450 19066
rect 4450 19014 4464 19066
rect 4488 19014 4502 19066
rect 4502 19014 4514 19066
rect 4514 19014 4544 19066
rect 4568 19014 4578 19066
rect 4578 19014 4624 19066
rect 4328 19012 4384 19014
rect 4408 19012 4464 19014
rect 4488 19012 4544 19014
rect 4568 19012 4624 19014
rect 3668 16346 3724 16348
rect 3748 16346 3804 16348
rect 3828 16346 3884 16348
rect 3908 16346 3964 16348
rect 3668 16294 3714 16346
rect 3714 16294 3724 16346
rect 3748 16294 3778 16346
rect 3778 16294 3790 16346
rect 3790 16294 3804 16346
rect 3828 16294 3842 16346
rect 3842 16294 3854 16346
rect 3854 16294 3884 16346
rect 3908 16294 3918 16346
rect 3918 16294 3964 16346
rect 3668 16292 3724 16294
rect 3748 16292 3804 16294
rect 3828 16292 3884 16294
rect 3908 16292 3964 16294
rect 4328 17978 4384 17980
rect 4408 17978 4464 17980
rect 4488 17978 4544 17980
rect 4568 17978 4624 17980
rect 4328 17926 4374 17978
rect 4374 17926 4384 17978
rect 4408 17926 4438 17978
rect 4438 17926 4450 17978
rect 4450 17926 4464 17978
rect 4488 17926 4502 17978
rect 4502 17926 4514 17978
rect 4514 17926 4544 17978
rect 4568 17926 4578 17978
rect 4578 17926 4624 17978
rect 4328 17924 4384 17926
rect 4408 17924 4464 17926
rect 4488 17924 4544 17926
rect 4568 17924 4624 17926
rect 4328 16890 4384 16892
rect 4408 16890 4464 16892
rect 4488 16890 4544 16892
rect 4568 16890 4624 16892
rect 4328 16838 4374 16890
rect 4374 16838 4384 16890
rect 4408 16838 4438 16890
rect 4438 16838 4450 16890
rect 4450 16838 4464 16890
rect 4488 16838 4502 16890
rect 4502 16838 4514 16890
rect 4514 16838 4544 16890
rect 4568 16838 4578 16890
rect 4578 16838 4624 16890
rect 4328 16836 4384 16838
rect 4408 16836 4464 16838
rect 4488 16836 4544 16838
rect 4568 16836 4624 16838
rect 3668 15258 3724 15260
rect 3748 15258 3804 15260
rect 3828 15258 3884 15260
rect 3908 15258 3964 15260
rect 3668 15206 3714 15258
rect 3714 15206 3724 15258
rect 3748 15206 3778 15258
rect 3778 15206 3790 15258
rect 3790 15206 3804 15258
rect 3828 15206 3842 15258
rect 3842 15206 3854 15258
rect 3854 15206 3884 15258
rect 3908 15206 3918 15258
rect 3918 15206 3964 15258
rect 3668 15204 3724 15206
rect 3748 15204 3804 15206
rect 3828 15204 3884 15206
rect 3908 15204 3964 15206
rect 4328 15802 4384 15804
rect 4408 15802 4464 15804
rect 4488 15802 4544 15804
rect 4568 15802 4624 15804
rect 4328 15750 4374 15802
rect 4374 15750 4384 15802
rect 4408 15750 4438 15802
rect 4438 15750 4450 15802
rect 4450 15750 4464 15802
rect 4488 15750 4502 15802
rect 4502 15750 4514 15802
rect 4514 15750 4544 15802
rect 4568 15750 4578 15802
rect 4578 15750 4624 15802
rect 4328 15748 4384 15750
rect 4408 15748 4464 15750
rect 4488 15748 4544 15750
rect 4568 15748 4624 15750
rect 4328 14714 4384 14716
rect 4408 14714 4464 14716
rect 4488 14714 4544 14716
rect 4568 14714 4624 14716
rect 4328 14662 4374 14714
rect 4374 14662 4384 14714
rect 4408 14662 4438 14714
rect 4438 14662 4450 14714
rect 4450 14662 4464 14714
rect 4488 14662 4502 14714
rect 4502 14662 4514 14714
rect 4514 14662 4544 14714
rect 4568 14662 4578 14714
rect 4578 14662 4624 14714
rect 4328 14660 4384 14662
rect 4408 14660 4464 14662
rect 4488 14660 4544 14662
rect 4568 14660 4624 14662
rect 3668 14170 3724 14172
rect 3748 14170 3804 14172
rect 3828 14170 3884 14172
rect 3908 14170 3964 14172
rect 3668 14118 3714 14170
rect 3714 14118 3724 14170
rect 3748 14118 3778 14170
rect 3778 14118 3790 14170
rect 3790 14118 3804 14170
rect 3828 14118 3842 14170
rect 3842 14118 3854 14170
rect 3854 14118 3884 14170
rect 3908 14118 3918 14170
rect 3918 14118 3964 14170
rect 3668 14116 3724 14118
rect 3748 14116 3804 14118
rect 3828 14116 3884 14118
rect 3908 14116 3964 14118
rect 4328 13626 4384 13628
rect 4408 13626 4464 13628
rect 4488 13626 4544 13628
rect 4568 13626 4624 13628
rect 4328 13574 4374 13626
rect 4374 13574 4384 13626
rect 4408 13574 4438 13626
rect 4438 13574 4450 13626
rect 4450 13574 4464 13626
rect 4488 13574 4502 13626
rect 4502 13574 4514 13626
rect 4514 13574 4544 13626
rect 4568 13574 4578 13626
rect 4578 13574 4624 13626
rect 4328 13572 4384 13574
rect 4408 13572 4464 13574
rect 4488 13572 4544 13574
rect 4568 13572 4624 13574
rect 3668 13082 3724 13084
rect 3748 13082 3804 13084
rect 3828 13082 3884 13084
rect 3908 13082 3964 13084
rect 3668 13030 3714 13082
rect 3714 13030 3724 13082
rect 3748 13030 3778 13082
rect 3778 13030 3790 13082
rect 3790 13030 3804 13082
rect 3828 13030 3842 13082
rect 3842 13030 3854 13082
rect 3854 13030 3884 13082
rect 3908 13030 3918 13082
rect 3918 13030 3964 13082
rect 3668 13028 3724 13030
rect 3748 13028 3804 13030
rect 3828 13028 3884 13030
rect 3908 13028 3964 13030
rect 4328 12538 4384 12540
rect 4408 12538 4464 12540
rect 4488 12538 4544 12540
rect 4568 12538 4624 12540
rect 4328 12486 4374 12538
rect 4374 12486 4384 12538
rect 4408 12486 4438 12538
rect 4438 12486 4450 12538
rect 4450 12486 4464 12538
rect 4488 12486 4502 12538
rect 4502 12486 4514 12538
rect 4514 12486 4544 12538
rect 4568 12486 4578 12538
rect 4578 12486 4624 12538
rect 4328 12484 4384 12486
rect 4408 12484 4464 12486
rect 4488 12484 4544 12486
rect 4568 12484 4624 12486
rect 5906 21292 5908 21312
rect 5908 21292 5960 21312
rect 5960 21292 5962 21312
rect 5906 21256 5962 21292
rect 3668 11994 3724 11996
rect 3748 11994 3804 11996
rect 3828 11994 3884 11996
rect 3908 11994 3964 11996
rect 3668 11942 3714 11994
rect 3714 11942 3724 11994
rect 3748 11942 3778 11994
rect 3778 11942 3790 11994
rect 3790 11942 3804 11994
rect 3828 11942 3842 11994
rect 3842 11942 3854 11994
rect 3854 11942 3884 11994
rect 3908 11942 3918 11994
rect 3918 11942 3964 11994
rect 3668 11940 3724 11942
rect 3748 11940 3804 11942
rect 3828 11940 3884 11942
rect 3908 11940 3964 11942
rect 4328 11450 4384 11452
rect 4408 11450 4464 11452
rect 4488 11450 4544 11452
rect 4568 11450 4624 11452
rect 4328 11398 4374 11450
rect 4374 11398 4384 11450
rect 4408 11398 4438 11450
rect 4438 11398 4450 11450
rect 4450 11398 4464 11450
rect 4488 11398 4502 11450
rect 4502 11398 4514 11450
rect 4514 11398 4544 11450
rect 4568 11398 4578 11450
rect 4578 11398 4624 11450
rect 4328 11396 4384 11398
rect 4408 11396 4464 11398
rect 4488 11396 4544 11398
rect 4568 11396 4624 11398
rect 3668 10906 3724 10908
rect 3748 10906 3804 10908
rect 3828 10906 3884 10908
rect 3908 10906 3964 10908
rect 3668 10854 3714 10906
rect 3714 10854 3724 10906
rect 3748 10854 3778 10906
rect 3778 10854 3790 10906
rect 3790 10854 3804 10906
rect 3828 10854 3842 10906
rect 3842 10854 3854 10906
rect 3854 10854 3884 10906
rect 3908 10854 3918 10906
rect 3918 10854 3964 10906
rect 3668 10852 3724 10854
rect 3748 10852 3804 10854
rect 3828 10852 3884 10854
rect 3908 10852 3964 10854
rect 4328 10362 4384 10364
rect 4408 10362 4464 10364
rect 4488 10362 4544 10364
rect 4568 10362 4624 10364
rect 4328 10310 4374 10362
rect 4374 10310 4384 10362
rect 4408 10310 4438 10362
rect 4438 10310 4450 10362
rect 4450 10310 4464 10362
rect 4488 10310 4502 10362
rect 4502 10310 4514 10362
rect 4514 10310 4544 10362
rect 4568 10310 4578 10362
rect 4578 10310 4624 10362
rect 4328 10308 4384 10310
rect 4408 10308 4464 10310
rect 4488 10308 4544 10310
rect 4568 10308 4624 10310
rect 3668 9818 3724 9820
rect 3748 9818 3804 9820
rect 3828 9818 3884 9820
rect 3908 9818 3964 9820
rect 3668 9766 3714 9818
rect 3714 9766 3724 9818
rect 3748 9766 3778 9818
rect 3778 9766 3790 9818
rect 3790 9766 3804 9818
rect 3828 9766 3842 9818
rect 3842 9766 3854 9818
rect 3854 9766 3884 9818
rect 3908 9766 3918 9818
rect 3918 9766 3964 9818
rect 3668 9764 3724 9766
rect 3748 9764 3804 9766
rect 3828 9764 3884 9766
rect 3908 9764 3964 9766
rect 4328 9274 4384 9276
rect 4408 9274 4464 9276
rect 4488 9274 4544 9276
rect 4568 9274 4624 9276
rect 4328 9222 4374 9274
rect 4374 9222 4384 9274
rect 4408 9222 4438 9274
rect 4438 9222 4450 9274
rect 4450 9222 4464 9274
rect 4488 9222 4502 9274
rect 4502 9222 4514 9274
rect 4514 9222 4544 9274
rect 4568 9222 4578 9274
rect 4578 9222 4624 9274
rect 4328 9220 4384 9222
rect 4408 9220 4464 9222
rect 4488 9220 4544 9222
rect 4568 9220 4624 9222
rect 3668 8730 3724 8732
rect 3748 8730 3804 8732
rect 3828 8730 3884 8732
rect 3908 8730 3964 8732
rect 3668 8678 3714 8730
rect 3714 8678 3724 8730
rect 3748 8678 3778 8730
rect 3778 8678 3790 8730
rect 3790 8678 3804 8730
rect 3828 8678 3842 8730
rect 3842 8678 3854 8730
rect 3854 8678 3884 8730
rect 3908 8678 3918 8730
rect 3918 8678 3964 8730
rect 3668 8676 3724 8678
rect 3748 8676 3804 8678
rect 3828 8676 3884 8678
rect 3908 8676 3964 8678
rect 7194 21936 7250 21992
rect 7286 21836 7288 21856
rect 7288 21836 7340 21856
rect 7340 21836 7342 21856
rect 7286 21800 7342 21836
rect 8574 21936 8630 21992
rect 10322 22380 10324 22400
rect 10324 22380 10376 22400
rect 10376 22380 10378 22400
rect 10322 22344 10378 22380
rect 9402 21256 9458 21312
rect 11702 21800 11758 21856
rect 4328 8186 4384 8188
rect 4408 8186 4464 8188
rect 4488 8186 4544 8188
rect 4568 8186 4624 8188
rect 4328 8134 4374 8186
rect 4374 8134 4384 8186
rect 4408 8134 4438 8186
rect 4438 8134 4450 8186
rect 4450 8134 4464 8186
rect 4488 8134 4502 8186
rect 4502 8134 4514 8186
rect 4514 8134 4544 8186
rect 4568 8134 4578 8186
rect 4578 8134 4624 8186
rect 4328 8132 4384 8134
rect 4408 8132 4464 8134
rect 4488 8132 4544 8134
rect 4568 8132 4624 8134
rect 3668 7642 3724 7644
rect 3748 7642 3804 7644
rect 3828 7642 3884 7644
rect 3908 7642 3964 7644
rect 3668 7590 3714 7642
rect 3714 7590 3724 7642
rect 3748 7590 3778 7642
rect 3778 7590 3790 7642
rect 3790 7590 3804 7642
rect 3828 7590 3842 7642
rect 3842 7590 3854 7642
rect 3854 7590 3884 7642
rect 3908 7590 3918 7642
rect 3918 7590 3964 7642
rect 3668 7588 3724 7590
rect 3748 7588 3804 7590
rect 3828 7588 3884 7590
rect 3908 7588 3964 7590
rect 3668 6554 3724 6556
rect 3748 6554 3804 6556
rect 3828 6554 3884 6556
rect 3908 6554 3964 6556
rect 3668 6502 3714 6554
rect 3714 6502 3724 6554
rect 3748 6502 3778 6554
rect 3778 6502 3790 6554
rect 3790 6502 3804 6554
rect 3828 6502 3842 6554
rect 3842 6502 3854 6554
rect 3854 6502 3884 6554
rect 3908 6502 3918 6554
rect 3918 6502 3964 6554
rect 3668 6500 3724 6502
rect 3748 6500 3804 6502
rect 3828 6500 3884 6502
rect 3908 6500 3964 6502
rect 4328 7098 4384 7100
rect 4408 7098 4464 7100
rect 4488 7098 4544 7100
rect 4568 7098 4624 7100
rect 4328 7046 4374 7098
rect 4374 7046 4384 7098
rect 4408 7046 4438 7098
rect 4438 7046 4450 7098
rect 4450 7046 4464 7098
rect 4488 7046 4502 7098
rect 4502 7046 4514 7098
rect 4514 7046 4544 7098
rect 4568 7046 4578 7098
rect 4578 7046 4624 7098
rect 4328 7044 4384 7046
rect 4408 7044 4464 7046
rect 4488 7044 4544 7046
rect 4568 7044 4624 7046
rect 4328 6010 4384 6012
rect 4408 6010 4464 6012
rect 4488 6010 4544 6012
rect 4568 6010 4624 6012
rect 4328 5958 4374 6010
rect 4374 5958 4384 6010
rect 4408 5958 4438 6010
rect 4438 5958 4450 6010
rect 4450 5958 4464 6010
rect 4488 5958 4502 6010
rect 4502 5958 4514 6010
rect 4514 5958 4544 6010
rect 4568 5958 4578 6010
rect 4578 5958 4624 6010
rect 4328 5956 4384 5958
rect 4408 5956 4464 5958
rect 4488 5956 4544 5958
rect 4568 5956 4624 5958
rect 3668 5466 3724 5468
rect 3748 5466 3804 5468
rect 3828 5466 3884 5468
rect 3908 5466 3964 5468
rect 3668 5414 3714 5466
rect 3714 5414 3724 5466
rect 3748 5414 3778 5466
rect 3778 5414 3790 5466
rect 3790 5414 3804 5466
rect 3828 5414 3842 5466
rect 3842 5414 3854 5466
rect 3854 5414 3884 5466
rect 3908 5414 3918 5466
rect 3918 5414 3964 5466
rect 3668 5412 3724 5414
rect 3748 5412 3804 5414
rect 3828 5412 3884 5414
rect 3908 5412 3964 5414
rect 14646 22344 14702 22400
rect 4328 4922 4384 4924
rect 4408 4922 4464 4924
rect 4488 4922 4544 4924
rect 4568 4922 4624 4924
rect 4328 4870 4374 4922
rect 4374 4870 4384 4922
rect 4408 4870 4438 4922
rect 4438 4870 4450 4922
rect 4450 4870 4464 4922
rect 4488 4870 4502 4922
rect 4502 4870 4514 4922
rect 4514 4870 4544 4922
rect 4568 4870 4578 4922
rect 4578 4870 4624 4922
rect 4328 4868 4384 4870
rect 4408 4868 4464 4870
rect 4488 4868 4544 4870
rect 4568 4868 4624 4870
rect 3668 4378 3724 4380
rect 3748 4378 3804 4380
rect 3828 4378 3884 4380
rect 3908 4378 3964 4380
rect 3668 4326 3714 4378
rect 3714 4326 3724 4378
rect 3748 4326 3778 4378
rect 3778 4326 3790 4378
rect 3790 4326 3804 4378
rect 3828 4326 3842 4378
rect 3842 4326 3854 4378
rect 3854 4326 3884 4378
rect 3908 4326 3918 4378
rect 3918 4326 3964 4378
rect 3668 4324 3724 4326
rect 3748 4324 3804 4326
rect 3828 4324 3884 4326
rect 3908 4324 3964 4326
rect 4328 3834 4384 3836
rect 4408 3834 4464 3836
rect 4488 3834 4544 3836
rect 4568 3834 4624 3836
rect 4328 3782 4374 3834
rect 4374 3782 4384 3834
rect 4408 3782 4438 3834
rect 4438 3782 4450 3834
rect 4450 3782 4464 3834
rect 4488 3782 4502 3834
rect 4502 3782 4514 3834
rect 4514 3782 4544 3834
rect 4568 3782 4578 3834
rect 4578 3782 4624 3834
rect 4328 3780 4384 3782
rect 4408 3780 4464 3782
rect 4488 3780 4544 3782
rect 4568 3780 4624 3782
rect 3668 3290 3724 3292
rect 3748 3290 3804 3292
rect 3828 3290 3884 3292
rect 3908 3290 3964 3292
rect 3668 3238 3714 3290
rect 3714 3238 3724 3290
rect 3748 3238 3778 3290
rect 3778 3238 3790 3290
rect 3790 3238 3804 3290
rect 3828 3238 3842 3290
rect 3842 3238 3854 3290
rect 3854 3238 3884 3290
rect 3908 3238 3918 3290
rect 3918 3238 3964 3290
rect 3668 3236 3724 3238
rect 3748 3236 3804 3238
rect 3828 3236 3884 3238
rect 3908 3236 3964 3238
rect 23018 19624 23074 19680
rect 23018 11736 23074 11792
rect 23018 3848 23074 3904
rect 4328 2746 4384 2748
rect 4408 2746 4464 2748
rect 4488 2746 4544 2748
rect 4568 2746 4624 2748
rect 4328 2694 4374 2746
rect 4374 2694 4384 2746
rect 4408 2694 4438 2746
rect 4438 2694 4450 2746
rect 4450 2694 4464 2746
rect 4488 2694 4502 2746
rect 4502 2694 4514 2746
rect 4514 2694 4544 2746
rect 4568 2694 4578 2746
rect 4578 2694 4624 2746
rect 4328 2692 4384 2694
rect 4408 2692 4464 2694
rect 4488 2692 4544 2694
rect 4568 2692 4624 2694
rect 3668 2202 3724 2204
rect 3748 2202 3804 2204
rect 3828 2202 3884 2204
rect 3908 2202 3964 2204
rect 3668 2150 3714 2202
rect 3714 2150 3724 2202
rect 3748 2150 3778 2202
rect 3778 2150 3790 2202
rect 3790 2150 3804 2202
rect 3828 2150 3842 2202
rect 3842 2150 3854 2202
rect 3854 2150 3884 2202
rect 3908 2150 3918 2202
rect 3918 2150 3964 2202
rect 3668 2148 3724 2150
rect 3748 2148 3804 2150
rect 3828 2148 3884 2150
rect 3908 2148 3964 2150
rect 4328 1658 4384 1660
rect 4408 1658 4464 1660
rect 4488 1658 4544 1660
rect 4568 1658 4624 1660
rect 4328 1606 4374 1658
rect 4374 1606 4384 1658
rect 4408 1606 4438 1658
rect 4438 1606 4450 1658
rect 4450 1606 4464 1658
rect 4488 1606 4502 1658
rect 4502 1606 4514 1658
rect 4514 1606 4544 1658
rect 4568 1606 4578 1658
rect 4578 1606 4624 1658
rect 4328 1604 4384 1606
rect 4408 1604 4464 1606
rect 4488 1604 4544 1606
rect 4568 1604 4624 1606
rect 3668 1114 3724 1116
rect 3748 1114 3804 1116
rect 3828 1114 3884 1116
rect 3908 1114 3964 1116
rect 3668 1062 3714 1114
rect 3714 1062 3724 1114
rect 3748 1062 3778 1114
rect 3778 1062 3790 1114
rect 3790 1062 3804 1114
rect 3828 1062 3842 1114
rect 3842 1062 3854 1114
rect 3854 1062 3884 1114
rect 3908 1062 3918 1114
rect 3918 1062 3964 1114
rect 3668 1060 3724 1062
rect 3748 1060 3804 1062
rect 3828 1060 3884 1062
rect 3908 1060 3964 1062
rect 4328 570 4384 572
rect 4408 570 4464 572
rect 4488 570 4544 572
rect 4568 570 4624 572
rect 4328 518 4374 570
rect 4374 518 4384 570
rect 4408 518 4438 570
rect 4438 518 4450 570
rect 4450 518 4464 570
rect 4488 518 4502 570
rect 4502 518 4514 570
rect 4514 518 4544 570
rect 4568 518 4578 570
rect 4578 518 4624 570
rect 4328 516 4384 518
rect 4408 516 4464 518
rect 4488 516 4544 518
rect 4568 516 4624 518
<< metal3 >>
rect 4318 23424 4634 23425
rect 4318 23360 4324 23424
rect 4388 23360 4404 23424
rect 4468 23360 4484 23424
rect 4548 23360 4564 23424
rect 4628 23360 4634 23424
rect 4318 23359 4634 23360
rect 3658 22880 3974 22881
rect 3658 22816 3664 22880
rect 3728 22816 3744 22880
rect 3808 22816 3824 22880
rect 3888 22816 3904 22880
rect 3968 22816 3974 22880
rect 3658 22815 3974 22816
rect 10317 22402 10383 22405
rect 14641 22402 14707 22405
rect 10317 22400 14707 22402
rect 10317 22344 10322 22400
rect 10378 22344 14646 22400
rect 14702 22344 14707 22400
rect 10317 22342 14707 22344
rect 10317 22339 10383 22342
rect 14641 22339 14707 22342
rect 4318 22336 4634 22337
rect 4318 22272 4324 22336
rect 4388 22272 4404 22336
rect 4468 22272 4484 22336
rect 4548 22272 4564 22336
rect 4628 22272 4634 22336
rect 4318 22271 4634 22272
rect 7189 21994 7255 21997
rect 8569 21994 8635 21997
rect 7189 21992 8635 21994
rect 7189 21936 7194 21992
rect 7250 21936 8574 21992
rect 8630 21936 8635 21992
rect 7189 21934 8635 21936
rect 7189 21931 7255 21934
rect 8569 21931 8635 21934
rect 7281 21858 7347 21861
rect 11697 21858 11763 21861
rect 7281 21856 11763 21858
rect 7281 21800 7286 21856
rect 7342 21800 11702 21856
rect 11758 21800 11763 21856
rect 7281 21798 11763 21800
rect 7281 21795 7347 21798
rect 11697 21795 11763 21798
rect 3658 21792 3974 21793
rect 3658 21728 3664 21792
rect 3728 21728 3744 21792
rect 3808 21728 3824 21792
rect 3888 21728 3904 21792
rect 3968 21728 3974 21792
rect 3658 21727 3974 21728
rect 5901 21314 5967 21317
rect 9397 21314 9463 21317
rect 5901 21312 9463 21314
rect 5901 21256 5906 21312
rect 5962 21256 9402 21312
rect 9458 21256 9463 21312
rect 5901 21254 9463 21256
rect 5901 21251 5967 21254
rect 9397 21251 9463 21254
rect 4318 21248 4634 21249
rect 4318 21184 4324 21248
rect 4388 21184 4404 21248
rect 4468 21184 4484 21248
rect 4548 21184 4564 21248
rect 4628 21184 4634 21248
rect 4318 21183 4634 21184
rect 3658 20704 3974 20705
rect 3658 20640 3664 20704
rect 3728 20640 3744 20704
rect 3808 20640 3824 20704
rect 3888 20640 3904 20704
rect 3968 20640 3974 20704
rect 3658 20639 3974 20640
rect 4318 20160 4634 20161
rect 4318 20096 4324 20160
rect 4388 20096 4404 20160
rect 4468 20096 4484 20160
rect 4548 20096 4564 20160
rect 4628 20096 4634 20160
rect 4318 20095 4634 20096
rect 23013 19682 23079 19685
rect 23600 19682 24000 19712
rect 23013 19680 24000 19682
rect 23013 19624 23018 19680
rect 23074 19624 24000 19680
rect 23013 19622 24000 19624
rect 23013 19619 23079 19622
rect 3658 19616 3974 19617
rect 3658 19552 3664 19616
rect 3728 19552 3744 19616
rect 3808 19552 3824 19616
rect 3888 19552 3904 19616
rect 3968 19552 3974 19616
rect 23600 19592 24000 19622
rect 3658 19551 3974 19552
rect 4318 19072 4634 19073
rect 4318 19008 4324 19072
rect 4388 19008 4404 19072
rect 4468 19008 4484 19072
rect 4548 19008 4564 19072
rect 4628 19008 4634 19072
rect 4318 19007 4634 19008
rect 3658 18528 3974 18529
rect 3658 18464 3664 18528
rect 3728 18464 3744 18528
rect 3808 18464 3824 18528
rect 3888 18464 3904 18528
rect 3968 18464 3974 18528
rect 3658 18463 3974 18464
rect 4318 17984 4634 17985
rect 4318 17920 4324 17984
rect 4388 17920 4404 17984
rect 4468 17920 4484 17984
rect 4548 17920 4564 17984
rect 4628 17920 4634 17984
rect 4318 17919 4634 17920
rect 3658 17440 3974 17441
rect 3658 17376 3664 17440
rect 3728 17376 3744 17440
rect 3808 17376 3824 17440
rect 3888 17376 3904 17440
rect 3968 17376 3974 17440
rect 3658 17375 3974 17376
rect 4318 16896 4634 16897
rect 4318 16832 4324 16896
rect 4388 16832 4404 16896
rect 4468 16832 4484 16896
rect 4548 16832 4564 16896
rect 4628 16832 4634 16896
rect 4318 16831 4634 16832
rect 3658 16352 3974 16353
rect 3658 16288 3664 16352
rect 3728 16288 3744 16352
rect 3808 16288 3824 16352
rect 3888 16288 3904 16352
rect 3968 16288 3974 16352
rect 3658 16287 3974 16288
rect 4318 15808 4634 15809
rect 4318 15744 4324 15808
rect 4388 15744 4404 15808
rect 4468 15744 4484 15808
rect 4548 15744 4564 15808
rect 4628 15744 4634 15808
rect 4318 15743 4634 15744
rect 3658 15264 3974 15265
rect 3658 15200 3664 15264
rect 3728 15200 3744 15264
rect 3808 15200 3824 15264
rect 3888 15200 3904 15264
rect 3968 15200 3974 15264
rect 3658 15199 3974 15200
rect 4318 14720 4634 14721
rect 4318 14656 4324 14720
rect 4388 14656 4404 14720
rect 4468 14656 4484 14720
rect 4548 14656 4564 14720
rect 4628 14656 4634 14720
rect 4318 14655 4634 14656
rect 3658 14176 3974 14177
rect 3658 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3904 14176
rect 3968 14112 3974 14176
rect 3658 14111 3974 14112
rect 4318 13632 4634 13633
rect 4318 13568 4324 13632
rect 4388 13568 4404 13632
rect 4468 13568 4484 13632
rect 4548 13568 4564 13632
rect 4628 13568 4634 13632
rect 4318 13567 4634 13568
rect 3658 13088 3974 13089
rect 3658 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3904 13088
rect 3968 13024 3974 13088
rect 3658 13023 3974 13024
rect 4318 12544 4634 12545
rect 4318 12480 4324 12544
rect 4388 12480 4404 12544
rect 4468 12480 4484 12544
rect 4548 12480 4564 12544
rect 4628 12480 4634 12544
rect 4318 12479 4634 12480
rect 3658 12000 3974 12001
rect 3658 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3904 12000
rect 3968 11936 3974 12000
rect 3658 11935 3974 11936
rect 23013 11794 23079 11797
rect 23600 11794 24000 11824
rect 23013 11792 24000 11794
rect 23013 11736 23018 11792
rect 23074 11736 24000 11792
rect 23013 11734 24000 11736
rect 23013 11731 23079 11734
rect 23600 11704 24000 11734
rect 4318 11456 4634 11457
rect 4318 11392 4324 11456
rect 4388 11392 4404 11456
rect 4468 11392 4484 11456
rect 4548 11392 4564 11456
rect 4628 11392 4634 11456
rect 4318 11391 4634 11392
rect 3658 10912 3974 10913
rect 3658 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3904 10912
rect 3968 10848 3974 10912
rect 3658 10847 3974 10848
rect 4318 10368 4634 10369
rect 4318 10304 4324 10368
rect 4388 10304 4404 10368
rect 4468 10304 4484 10368
rect 4548 10304 4564 10368
rect 4628 10304 4634 10368
rect 4318 10303 4634 10304
rect 3658 9824 3974 9825
rect 3658 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3904 9824
rect 3968 9760 3974 9824
rect 3658 9759 3974 9760
rect 4318 9280 4634 9281
rect 4318 9216 4324 9280
rect 4388 9216 4404 9280
rect 4468 9216 4484 9280
rect 4548 9216 4564 9280
rect 4628 9216 4634 9280
rect 4318 9215 4634 9216
rect 3658 8736 3974 8737
rect 3658 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3904 8736
rect 3968 8672 3974 8736
rect 3658 8671 3974 8672
rect 4318 8192 4634 8193
rect 4318 8128 4324 8192
rect 4388 8128 4404 8192
rect 4468 8128 4484 8192
rect 4548 8128 4564 8192
rect 4628 8128 4634 8192
rect 4318 8127 4634 8128
rect 3658 7648 3974 7649
rect 3658 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3904 7648
rect 3968 7584 3974 7648
rect 3658 7583 3974 7584
rect 4318 7104 4634 7105
rect 4318 7040 4324 7104
rect 4388 7040 4404 7104
rect 4468 7040 4484 7104
rect 4548 7040 4564 7104
rect 4628 7040 4634 7104
rect 4318 7039 4634 7040
rect 3658 6560 3974 6561
rect 3658 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3974 6560
rect 3658 6495 3974 6496
rect 4318 6016 4634 6017
rect 4318 5952 4324 6016
rect 4388 5952 4404 6016
rect 4468 5952 4484 6016
rect 4548 5952 4564 6016
rect 4628 5952 4634 6016
rect 4318 5951 4634 5952
rect 3658 5472 3974 5473
rect 3658 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3974 5472
rect 3658 5407 3974 5408
rect 4318 4928 4634 4929
rect 4318 4864 4324 4928
rect 4388 4864 4404 4928
rect 4468 4864 4484 4928
rect 4548 4864 4564 4928
rect 4628 4864 4634 4928
rect 4318 4863 4634 4864
rect 3658 4384 3974 4385
rect 3658 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3974 4384
rect 3658 4319 3974 4320
rect 23013 3906 23079 3909
rect 23600 3906 24000 3936
rect 23013 3904 24000 3906
rect 23013 3848 23018 3904
rect 23074 3848 24000 3904
rect 23013 3846 24000 3848
rect 23013 3843 23079 3846
rect 4318 3840 4634 3841
rect 4318 3776 4324 3840
rect 4388 3776 4404 3840
rect 4468 3776 4484 3840
rect 4548 3776 4564 3840
rect 4628 3776 4634 3840
rect 23600 3816 24000 3846
rect 4318 3775 4634 3776
rect 3658 3296 3974 3297
rect 3658 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3974 3296
rect 3658 3231 3974 3232
rect 4318 2752 4634 2753
rect 4318 2688 4324 2752
rect 4388 2688 4404 2752
rect 4468 2688 4484 2752
rect 4548 2688 4564 2752
rect 4628 2688 4634 2752
rect 4318 2687 4634 2688
rect 3658 2208 3974 2209
rect 3658 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3974 2208
rect 3658 2143 3974 2144
rect 4318 1664 4634 1665
rect 4318 1600 4324 1664
rect 4388 1600 4404 1664
rect 4468 1600 4484 1664
rect 4548 1600 4564 1664
rect 4628 1600 4634 1664
rect 4318 1599 4634 1600
rect 3658 1120 3974 1121
rect 3658 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3974 1120
rect 3658 1055 3974 1056
rect 4318 576 4634 577
rect 4318 512 4324 576
rect 4388 512 4404 576
rect 4468 512 4484 576
rect 4548 512 4564 576
rect 4628 512 4634 576
rect 4318 511 4634 512
<< via3 >>
rect 4324 23420 4388 23424
rect 4324 23364 4328 23420
rect 4328 23364 4384 23420
rect 4384 23364 4388 23420
rect 4324 23360 4388 23364
rect 4404 23420 4468 23424
rect 4404 23364 4408 23420
rect 4408 23364 4464 23420
rect 4464 23364 4468 23420
rect 4404 23360 4468 23364
rect 4484 23420 4548 23424
rect 4484 23364 4488 23420
rect 4488 23364 4544 23420
rect 4544 23364 4548 23420
rect 4484 23360 4548 23364
rect 4564 23420 4628 23424
rect 4564 23364 4568 23420
rect 4568 23364 4624 23420
rect 4624 23364 4628 23420
rect 4564 23360 4628 23364
rect 3664 22876 3728 22880
rect 3664 22820 3668 22876
rect 3668 22820 3724 22876
rect 3724 22820 3728 22876
rect 3664 22816 3728 22820
rect 3744 22876 3808 22880
rect 3744 22820 3748 22876
rect 3748 22820 3804 22876
rect 3804 22820 3808 22876
rect 3744 22816 3808 22820
rect 3824 22876 3888 22880
rect 3824 22820 3828 22876
rect 3828 22820 3884 22876
rect 3884 22820 3888 22876
rect 3824 22816 3888 22820
rect 3904 22876 3968 22880
rect 3904 22820 3908 22876
rect 3908 22820 3964 22876
rect 3964 22820 3968 22876
rect 3904 22816 3968 22820
rect 4324 22332 4388 22336
rect 4324 22276 4328 22332
rect 4328 22276 4384 22332
rect 4384 22276 4388 22332
rect 4324 22272 4388 22276
rect 4404 22332 4468 22336
rect 4404 22276 4408 22332
rect 4408 22276 4464 22332
rect 4464 22276 4468 22332
rect 4404 22272 4468 22276
rect 4484 22332 4548 22336
rect 4484 22276 4488 22332
rect 4488 22276 4544 22332
rect 4544 22276 4548 22332
rect 4484 22272 4548 22276
rect 4564 22332 4628 22336
rect 4564 22276 4568 22332
rect 4568 22276 4624 22332
rect 4624 22276 4628 22332
rect 4564 22272 4628 22276
rect 3664 21788 3728 21792
rect 3664 21732 3668 21788
rect 3668 21732 3724 21788
rect 3724 21732 3728 21788
rect 3664 21728 3728 21732
rect 3744 21788 3808 21792
rect 3744 21732 3748 21788
rect 3748 21732 3804 21788
rect 3804 21732 3808 21788
rect 3744 21728 3808 21732
rect 3824 21788 3888 21792
rect 3824 21732 3828 21788
rect 3828 21732 3884 21788
rect 3884 21732 3888 21788
rect 3824 21728 3888 21732
rect 3904 21788 3968 21792
rect 3904 21732 3908 21788
rect 3908 21732 3964 21788
rect 3964 21732 3968 21788
rect 3904 21728 3968 21732
rect 4324 21244 4388 21248
rect 4324 21188 4328 21244
rect 4328 21188 4384 21244
rect 4384 21188 4388 21244
rect 4324 21184 4388 21188
rect 4404 21244 4468 21248
rect 4404 21188 4408 21244
rect 4408 21188 4464 21244
rect 4464 21188 4468 21244
rect 4404 21184 4468 21188
rect 4484 21244 4548 21248
rect 4484 21188 4488 21244
rect 4488 21188 4544 21244
rect 4544 21188 4548 21244
rect 4484 21184 4548 21188
rect 4564 21244 4628 21248
rect 4564 21188 4568 21244
rect 4568 21188 4624 21244
rect 4624 21188 4628 21244
rect 4564 21184 4628 21188
rect 3664 20700 3728 20704
rect 3664 20644 3668 20700
rect 3668 20644 3724 20700
rect 3724 20644 3728 20700
rect 3664 20640 3728 20644
rect 3744 20700 3808 20704
rect 3744 20644 3748 20700
rect 3748 20644 3804 20700
rect 3804 20644 3808 20700
rect 3744 20640 3808 20644
rect 3824 20700 3888 20704
rect 3824 20644 3828 20700
rect 3828 20644 3884 20700
rect 3884 20644 3888 20700
rect 3824 20640 3888 20644
rect 3904 20700 3968 20704
rect 3904 20644 3908 20700
rect 3908 20644 3964 20700
rect 3964 20644 3968 20700
rect 3904 20640 3968 20644
rect 4324 20156 4388 20160
rect 4324 20100 4328 20156
rect 4328 20100 4384 20156
rect 4384 20100 4388 20156
rect 4324 20096 4388 20100
rect 4404 20156 4468 20160
rect 4404 20100 4408 20156
rect 4408 20100 4464 20156
rect 4464 20100 4468 20156
rect 4404 20096 4468 20100
rect 4484 20156 4548 20160
rect 4484 20100 4488 20156
rect 4488 20100 4544 20156
rect 4544 20100 4548 20156
rect 4484 20096 4548 20100
rect 4564 20156 4628 20160
rect 4564 20100 4568 20156
rect 4568 20100 4624 20156
rect 4624 20100 4628 20156
rect 4564 20096 4628 20100
rect 3664 19612 3728 19616
rect 3664 19556 3668 19612
rect 3668 19556 3724 19612
rect 3724 19556 3728 19612
rect 3664 19552 3728 19556
rect 3744 19612 3808 19616
rect 3744 19556 3748 19612
rect 3748 19556 3804 19612
rect 3804 19556 3808 19612
rect 3744 19552 3808 19556
rect 3824 19612 3888 19616
rect 3824 19556 3828 19612
rect 3828 19556 3884 19612
rect 3884 19556 3888 19612
rect 3824 19552 3888 19556
rect 3904 19612 3968 19616
rect 3904 19556 3908 19612
rect 3908 19556 3964 19612
rect 3964 19556 3968 19612
rect 3904 19552 3968 19556
rect 4324 19068 4388 19072
rect 4324 19012 4328 19068
rect 4328 19012 4384 19068
rect 4384 19012 4388 19068
rect 4324 19008 4388 19012
rect 4404 19068 4468 19072
rect 4404 19012 4408 19068
rect 4408 19012 4464 19068
rect 4464 19012 4468 19068
rect 4404 19008 4468 19012
rect 4484 19068 4548 19072
rect 4484 19012 4488 19068
rect 4488 19012 4544 19068
rect 4544 19012 4548 19068
rect 4484 19008 4548 19012
rect 4564 19068 4628 19072
rect 4564 19012 4568 19068
rect 4568 19012 4624 19068
rect 4624 19012 4628 19068
rect 4564 19008 4628 19012
rect 3664 18524 3728 18528
rect 3664 18468 3668 18524
rect 3668 18468 3724 18524
rect 3724 18468 3728 18524
rect 3664 18464 3728 18468
rect 3744 18524 3808 18528
rect 3744 18468 3748 18524
rect 3748 18468 3804 18524
rect 3804 18468 3808 18524
rect 3744 18464 3808 18468
rect 3824 18524 3888 18528
rect 3824 18468 3828 18524
rect 3828 18468 3884 18524
rect 3884 18468 3888 18524
rect 3824 18464 3888 18468
rect 3904 18524 3968 18528
rect 3904 18468 3908 18524
rect 3908 18468 3964 18524
rect 3964 18468 3968 18524
rect 3904 18464 3968 18468
rect 4324 17980 4388 17984
rect 4324 17924 4328 17980
rect 4328 17924 4384 17980
rect 4384 17924 4388 17980
rect 4324 17920 4388 17924
rect 4404 17980 4468 17984
rect 4404 17924 4408 17980
rect 4408 17924 4464 17980
rect 4464 17924 4468 17980
rect 4404 17920 4468 17924
rect 4484 17980 4548 17984
rect 4484 17924 4488 17980
rect 4488 17924 4544 17980
rect 4544 17924 4548 17980
rect 4484 17920 4548 17924
rect 4564 17980 4628 17984
rect 4564 17924 4568 17980
rect 4568 17924 4624 17980
rect 4624 17924 4628 17980
rect 4564 17920 4628 17924
rect 3664 17436 3728 17440
rect 3664 17380 3668 17436
rect 3668 17380 3724 17436
rect 3724 17380 3728 17436
rect 3664 17376 3728 17380
rect 3744 17436 3808 17440
rect 3744 17380 3748 17436
rect 3748 17380 3804 17436
rect 3804 17380 3808 17436
rect 3744 17376 3808 17380
rect 3824 17436 3888 17440
rect 3824 17380 3828 17436
rect 3828 17380 3884 17436
rect 3884 17380 3888 17436
rect 3824 17376 3888 17380
rect 3904 17436 3968 17440
rect 3904 17380 3908 17436
rect 3908 17380 3964 17436
rect 3964 17380 3968 17436
rect 3904 17376 3968 17380
rect 4324 16892 4388 16896
rect 4324 16836 4328 16892
rect 4328 16836 4384 16892
rect 4384 16836 4388 16892
rect 4324 16832 4388 16836
rect 4404 16892 4468 16896
rect 4404 16836 4408 16892
rect 4408 16836 4464 16892
rect 4464 16836 4468 16892
rect 4404 16832 4468 16836
rect 4484 16892 4548 16896
rect 4484 16836 4488 16892
rect 4488 16836 4544 16892
rect 4544 16836 4548 16892
rect 4484 16832 4548 16836
rect 4564 16892 4628 16896
rect 4564 16836 4568 16892
rect 4568 16836 4624 16892
rect 4624 16836 4628 16892
rect 4564 16832 4628 16836
rect 3664 16348 3728 16352
rect 3664 16292 3668 16348
rect 3668 16292 3724 16348
rect 3724 16292 3728 16348
rect 3664 16288 3728 16292
rect 3744 16348 3808 16352
rect 3744 16292 3748 16348
rect 3748 16292 3804 16348
rect 3804 16292 3808 16348
rect 3744 16288 3808 16292
rect 3824 16348 3888 16352
rect 3824 16292 3828 16348
rect 3828 16292 3884 16348
rect 3884 16292 3888 16348
rect 3824 16288 3888 16292
rect 3904 16348 3968 16352
rect 3904 16292 3908 16348
rect 3908 16292 3964 16348
rect 3964 16292 3968 16348
rect 3904 16288 3968 16292
rect 4324 15804 4388 15808
rect 4324 15748 4328 15804
rect 4328 15748 4384 15804
rect 4384 15748 4388 15804
rect 4324 15744 4388 15748
rect 4404 15804 4468 15808
rect 4404 15748 4408 15804
rect 4408 15748 4464 15804
rect 4464 15748 4468 15804
rect 4404 15744 4468 15748
rect 4484 15804 4548 15808
rect 4484 15748 4488 15804
rect 4488 15748 4544 15804
rect 4544 15748 4548 15804
rect 4484 15744 4548 15748
rect 4564 15804 4628 15808
rect 4564 15748 4568 15804
rect 4568 15748 4624 15804
rect 4624 15748 4628 15804
rect 4564 15744 4628 15748
rect 3664 15260 3728 15264
rect 3664 15204 3668 15260
rect 3668 15204 3724 15260
rect 3724 15204 3728 15260
rect 3664 15200 3728 15204
rect 3744 15260 3808 15264
rect 3744 15204 3748 15260
rect 3748 15204 3804 15260
rect 3804 15204 3808 15260
rect 3744 15200 3808 15204
rect 3824 15260 3888 15264
rect 3824 15204 3828 15260
rect 3828 15204 3884 15260
rect 3884 15204 3888 15260
rect 3824 15200 3888 15204
rect 3904 15260 3968 15264
rect 3904 15204 3908 15260
rect 3908 15204 3964 15260
rect 3964 15204 3968 15260
rect 3904 15200 3968 15204
rect 4324 14716 4388 14720
rect 4324 14660 4328 14716
rect 4328 14660 4384 14716
rect 4384 14660 4388 14716
rect 4324 14656 4388 14660
rect 4404 14716 4468 14720
rect 4404 14660 4408 14716
rect 4408 14660 4464 14716
rect 4464 14660 4468 14716
rect 4404 14656 4468 14660
rect 4484 14716 4548 14720
rect 4484 14660 4488 14716
rect 4488 14660 4544 14716
rect 4544 14660 4548 14716
rect 4484 14656 4548 14660
rect 4564 14716 4628 14720
rect 4564 14660 4568 14716
rect 4568 14660 4624 14716
rect 4624 14660 4628 14716
rect 4564 14656 4628 14660
rect 3664 14172 3728 14176
rect 3664 14116 3668 14172
rect 3668 14116 3724 14172
rect 3724 14116 3728 14172
rect 3664 14112 3728 14116
rect 3744 14172 3808 14176
rect 3744 14116 3748 14172
rect 3748 14116 3804 14172
rect 3804 14116 3808 14172
rect 3744 14112 3808 14116
rect 3824 14172 3888 14176
rect 3824 14116 3828 14172
rect 3828 14116 3884 14172
rect 3884 14116 3888 14172
rect 3824 14112 3888 14116
rect 3904 14172 3968 14176
rect 3904 14116 3908 14172
rect 3908 14116 3964 14172
rect 3964 14116 3968 14172
rect 3904 14112 3968 14116
rect 4324 13628 4388 13632
rect 4324 13572 4328 13628
rect 4328 13572 4384 13628
rect 4384 13572 4388 13628
rect 4324 13568 4388 13572
rect 4404 13628 4468 13632
rect 4404 13572 4408 13628
rect 4408 13572 4464 13628
rect 4464 13572 4468 13628
rect 4404 13568 4468 13572
rect 4484 13628 4548 13632
rect 4484 13572 4488 13628
rect 4488 13572 4544 13628
rect 4544 13572 4548 13628
rect 4484 13568 4548 13572
rect 4564 13628 4628 13632
rect 4564 13572 4568 13628
rect 4568 13572 4624 13628
rect 4624 13572 4628 13628
rect 4564 13568 4628 13572
rect 3664 13084 3728 13088
rect 3664 13028 3668 13084
rect 3668 13028 3724 13084
rect 3724 13028 3728 13084
rect 3664 13024 3728 13028
rect 3744 13084 3808 13088
rect 3744 13028 3748 13084
rect 3748 13028 3804 13084
rect 3804 13028 3808 13084
rect 3744 13024 3808 13028
rect 3824 13084 3888 13088
rect 3824 13028 3828 13084
rect 3828 13028 3884 13084
rect 3884 13028 3888 13084
rect 3824 13024 3888 13028
rect 3904 13084 3968 13088
rect 3904 13028 3908 13084
rect 3908 13028 3964 13084
rect 3964 13028 3968 13084
rect 3904 13024 3968 13028
rect 4324 12540 4388 12544
rect 4324 12484 4328 12540
rect 4328 12484 4384 12540
rect 4384 12484 4388 12540
rect 4324 12480 4388 12484
rect 4404 12540 4468 12544
rect 4404 12484 4408 12540
rect 4408 12484 4464 12540
rect 4464 12484 4468 12540
rect 4404 12480 4468 12484
rect 4484 12540 4548 12544
rect 4484 12484 4488 12540
rect 4488 12484 4544 12540
rect 4544 12484 4548 12540
rect 4484 12480 4548 12484
rect 4564 12540 4628 12544
rect 4564 12484 4568 12540
rect 4568 12484 4624 12540
rect 4624 12484 4628 12540
rect 4564 12480 4628 12484
rect 3664 11996 3728 12000
rect 3664 11940 3668 11996
rect 3668 11940 3724 11996
rect 3724 11940 3728 11996
rect 3664 11936 3728 11940
rect 3744 11996 3808 12000
rect 3744 11940 3748 11996
rect 3748 11940 3804 11996
rect 3804 11940 3808 11996
rect 3744 11936 3808 11940
rect 3824 11996 3888 12000
rect 3824 11940 3828 11996
rect 3828 11940 3884 11996
rect 3884 11940 3888 11996
rect 3824 11936 3888 11940
rect 3904 11996 3968 12000
rect 3904 11940 3908 11996
rect 3908 11940 3964 11996
rect 3964 11940 3968 11996
rect 3904 11936 3968 11940
rect 4324 11452 4388 11456
rect 4324 11396 4328 11452
rect 4328 11396 4384 11452
rect 4384 11396 4388 11452
rect 4324 11392 4388 11396
rect 4404 11452 4468 11456
rect 4404 11396 4408 11452
rect 4408 11396 4464 11452
rect 4464 11396 4468 11452
rect 4404 11392 4468 11396
rect 4484 11452 4548 11456
rect 4484 11396 4488 11452
rect 4488 11396 4544 11452
rect 4544 11396 4548 11452
rect 4484 11392 4548 11396
rect 4564 11452 4628 11456
rect 4564 11396 4568 11452
rect 4568 11396 4624 11452
rect 4624 11396 4628 11452
rect 4564 11392 4628 11396
rect 3664 10908 3728 10912
rect 3664 10852 3668 10908
rect 3668 10852 3724 10908
rect 3724 10852 3728 10908
rect 3664 10848 3728 10852
rect 3744 10908 3808 10912
rect 3744 10852 3748 10908
rect 3748 10852 3804 10908
rect 3804 10852 3808 10908
rect 3744 10848 3808 10852
rect 3824 10908 3888 10912
rect 3824 10852 3828 10908
rect 3828 10852 3884 10908
rect 3884 10852 3888 10908
rect 3824 10848 3888 10852
rect 3904 10908 3968 10912
rect 3904 10852 3908 10908
rect 3908 10852 3964 10908
rect 3964 10852 3968 10908
rect 3904 10848 3968 10852
rect 4324 10364 4388 10368
rect 4324 10308 4328 10364
rect 4328 10308 4384 10364
rect 4384 10308 4388 10364
rect 4324 10304 4388 10308
rect 4404 10364 4468 10368
rect 4404 10308 4408 10364
rect 4408 10308 4464 10364
rect 4464 10308 4468 10364
rect 4404 10304 4468 10308
rect 4484 10364 4548 10368
rect 4484 10308 4488 10364
rect 4488 10308 4544 10364
rect 4544 10308 4548 10364
rect 4484 10304 4548 10308
rect 4564 10364 4628 10368
rect 4564 10308 4568 10364
rect 4568 10308 4624 10364
rect 4624 10308 4628 10364
rect 4564 10304 4628 10308
rect 3664 9820 3728 9824
rect 3664 9764 3668 9820
rect 3668 9764 3724 9820
rect 3724 9764 3728 9820
rect 3664 9760 3728 9764
rect 3744 9820 3808 9824
rect 3744 9764 3748 9820
rect 3748 9764 3804 9820
rect 3804 9764 3808 9820
rect 3744 9760 3808 9764
rect 3824 9820 3888 9824
rect 3824 9764 3828 9820
rect 3828 9764 3884 9820
rect 3884 9764 3888 9820
rect 3824 9760 3888 9764
rect 3904 9820 3968 9824
rect 3904 9764 3908 9820
rect 3908 9764 3964 9820
rect 3964 9764 3968 9820
rect 3904 9760 3968 9764
rect 4324 9276 4388 9280
rect 4324 9220 4328 9276
rect 4328 9220 4384 9276
rect 4384 9220 4388 9276
rect 4324 9216 4388 9220
rect 4404 9276 4468 9280
rect 4404 9220 4408 9276
rect 4408 9220 4464 9276
rect 4464 9220 4468 9276
rect 4404 9216 4468 9220
rect 4484 9276 4548 9280
rect 4484 9220 4488 9276
rect 4488 9220 4544 9276
rect 4544 9220 4548 9276
rect 4484 9216 4548 9220
rect 4564 9276 4628 9280
rect 4564 9220 4568 9276
rect 4568 9220 4624 9276
rect 4624 9220 4628 9276
rect 4564 9216 4628 9220
rect 3664 8732 3728 8736
rect 3664 8676 3668 8732
rect 3668 8676 3724 8732
rect 3724 8676 3728 8732
rect 3664 8672 3728 8676
rect 3744 8732 3808 8736
rect 3744 8676 3748 8732
rect 3748 8676 3804 8732
rect 3804 8676 3808 8732
rect 3744 8672 3808 8676
rect 3824 8732 3888 8736
rect 3824 8676 3828 8732
rect 3828 8676 3884 8732
rect 3884 8676 3888 8732
rect 3824 8672 3888 8676
rect 3904 8732 3968 8736
rect 3904 8676 3908 8732
rect 3908 8676 3964 8732
rect 3964 8676 3968 8732
rect 3904 8672 3968 8676
rect 4324 8188 4388 8192
rect 4324 8132 4328 8188
rect 4328 8132 4384 8188
rect 4384 8132 4388 8188
rect 4324 8128 4388 8132
rect 4404 8188 4468 8192
rect 4404 8132 4408 8188
rect 4408 8132 4464 8188
rect 4464 8132 4468 8188
rect 4404 8128 4468 8132
rect 4484 8188 4548 8192
rect 4484 8132 4488 8188
rect 4488 8132 4544 8188
rect 4544 8132 4548 8188
rect 4484 8128 4548 8132
rect 4564 8188 4628 8192
rect 4564 8132 4568 8188
rect 4568 8132 4624 8188
rect 4624 8132 4628 8188
rect 4564 8128 4628 8132
rect 3664 7644 3728 7648
rect 3664 7588 3668 7644
rect 3668 7588 3724 7644
rect 3724 7588 3728 7644
rect 3664 7584 3728 7588
rect 3744 7644 3808 7648
rect 3744 7588 3748 7644
rect 3748 7588 3804 7644
rect 3804 7588 3808 7644
rect 3744 7584 3808 7588
rect 3824 7644 3888 7648
rect 3824 7588 3828 7644
rect 3828 7588 3884 7644
rect 3884 7588 3888 7644
rect 3824 7584 3888 7588
rect 3904 7644 3968 7648
rect 3904 7588 3908 7644
rect 3908 7588 3964 7644
rect 3964 7588 3968 7644
rect 3904 7584 3968 7588
rect 4324 7100 4388 7104
rect 4324 7044 4328 7100
rect 4328 7044 4384 7100
rect 4384 7044 4388 7100
rect 4324 7040 4388 7044
rect 4404 7100 4468 7104
rect 4404 7044 4408 7100
rect 4408 7044 4464 7100
rect 4464 7044 4468 7100
rect 4404 7040 4468 7044
rect 4484 7100 4548 7104
rect 4484 7044 4488 7100
rect 4488 7044 4544 7100
rect 4544 7044 4548 7100
rect 4484 7040 4548 7044
rect 4564 7100 4628 7104
rect 4564 7044 4568 7100
rect 4568 7044 4624 7100
rect 4624 7044 4628 7100
rect 4564 7040 4628 7044
rect 3664 6556 3728 6560
rect 3664 6500 3668 6556
rect 3668 6500 3724 6556
rect 3724 6500 3728 6556
rect 3664 6496 3728 6500
rect 3744 6556 3808 6560
rect 3744 6500 3748 6556
rect 3748 6500 3804 6556
rect 3804 6500 3808 6556
rect 3744 6496 3808 6500
rect 3824 6556 3888 6560
rect 3824 6500 3828 6556
rect 3828 6500 3884 6556
rect 3884 6500 3888 6556
rect 3824 6496 3888 6500
rect 3904 6556 3968 6560
rect 3904 6500 3908 6556
rect 3908 6500 3964 6556
rect 3964 6500 3968 6556
rect 3904 6496 3968 6500
rect 4324 6012 4388 6016
rect 4324 5956 4328 6012
rect 4328 5956 4384 6012
rect 4384 5956 4388 6012
rect 4324 5952 4388 5956
rect 4404 6012 4468 6016
rect 4404 5956 4408 6012
rect 4408 5956 4464 6012
rect 4464 5956 4468 6012
rect 4404 5952 4468 5956
rect 4484 6012 4548 6016
rect 4484 5956 4488 6012
rect 4488 5956 4544 6012
rect 4544 5956 4548 6012
rect 4484 5952 4548 5956
rect 4564 6012 4628 6016
rect 4564 5956 4568 6012
rect 4568 5956 4624 6012
rect 4624 5956 4628 6012
rect 4564 5952 4628 5956
rect 3664 5468 3728 5472
rect 3664 5412 3668 5468
rect 3668 5412 3724 5468
rect 3724 5412 3728 5468
rect 3664 5408 3728 5412
rect 3744 5468 3808 5472
rect 3744 5412 3748 5468
rect 3748 5412 3804 5468
rect 3804 5412 3808 5468
rect 3744 5408 3808 5412
rect 3824 5468 3888 5472
rect 3824 5412 3828 5468
rect 3828 5412 3884 5468
rect 3884 5412 3888 5468
rect 3824 5408 3888 5412
rect 3904 5468 3968 5472
rect 3904 5412 3908 5468
rect 3908 5412 3964 5468
rect 3964 5412 3968 5468
rect 3904 5408 3968 5412
rect 4324 4924 4388 4928
rect 4324 4868 4328 4924
rect 4328 4868 4384 4924
rect 4384 4868 4388 4924
rect 4324 4864 4388 4868
rect 4404 4924 4468 4928
rect 4404 4868 4408 4924
rect 4408 4868 4464 4924
rect 4464 4868 4468 4924
rect 4404 4864 4468 4868
rect 4484 4924 4548 4928
rect 4484 4868 4488 4924
rect 4488 4868 4544 4924
rect 4544 4868 4548 4924
rect 4484 4864 4548 4868
rect 4564 4924 4628 4928
rect 4564 4868 4568 4924
rect 4568 4868 4624 4924
rect 4624 4868 4628 4924
rect 4564 4864 4628 4868
rect 3664 4380 3728 4384
rect 3664 4324 3668 4380
rect 3668 4324 3724 4380
rect 3724 4324 3728 4380
rect 3664 4320 3728 4324
rect 3744 4380 3808 4384
rect 3744 4324 3748 4380
rect 3748 4324 3804 4380
rect 3804 4324 3808 4380
rect 3744 4320 3808 4324
rect 3824 4380 3888 4384
rect 3824 4324 3828 4380
rect 3828 4324 3884 4380
rect 3884 4324 3888 4380
rect 3824 4320 3888 4324
rect 3904 4380 3968 4384
rect 3904 4324 3908 4380
rect 3908 4324 3964 4380
rect 3964 4324 3968 4380
rect 3904 4320 3968 4324
rect 4324 3836 4388 3840
rect 4324 3780 4328 3836
rect 4328 3780 4384 3836
rect 4384 3780 4388 3836
rect 4324 3776 4388 3780
rect 4404 3836 4468 3840
rect 4404 3780 4408 3836
rect 4408 3780 4464 3836
rect 4464 3780 4468 3836
rect 4404 3776 4468 3780
rect 4484 3836 4548 3840
rect 4484 3780 4488 3836
rect 4488 3780 4544 3836
rect 4544 3780 4548 3836
rect 4484 3776 4548 3780
rect 4564 3836 4628 3840
rect 4564 3780 4568 3836
rect 4568 3780 4624 3836
rect 4624 3780 4628 3836
rect 4564 3776 4628 3780
rect 3664 3292 3728 3296
rect 3664 3236 3668 3292
rect 3668 3236 3724 3292
rect 3724 3236 3728 3292
rect 3664 3232 3728 3236
rect 3744 3292 3808 3296
rect 3744 3236 3748 3292
rect 3748 3236 3804 3292
rect 3804 3236 3808 3292
rect 3744 3232 3808 3236
rect 3824 3292 3888 3296
rect 3824 3236 3828 3292
rect 3828 3236 3884 3292
rect 3884 3236 3888 3292
rect 3824 3232 3888 3236
rect 3904 3292 3968 3296
rect 3904 3236 3908 3292
rect 3908 3236 3964 3292
rect 3964 3236 3968 3292
rect 3904 3232 3968 3236
rect 4324 2748 4388 2752
rect 4324 2692 4328 2748
rect 4328 2692 4384 2748
rect 4384 2692 4388 2748
rect 4324 2688 4388 2692
rect 4404 2748 4468 2752
rect 4404 2692 4408 2748
rect 4408 2692 4464 2748
rect 4464 2692 4468 2748
rect 4404 2688 4468 2692
rect 4484 2748 4548 2752
rect 4484 2692 4488 2748
rect 4488 2692 4544 2748
rect 4544 2692 4548 2748
rect 4484 2688 4548 2692
rect 4564 2748 4628 2752
rect 4564 2692 4568 2748
rect 4568 2692 4624 2748
rect 4624 2692 4628 2748
rect 4564 2688 4628 2692
rect 3664 2204 3728 2208
rect 3664 2148 3668 2204
rect 3668 2148 3724 2204
rect 3724 2148 3728 2204
rect 3664 2144 3728 2148
rect 3744 2204 3808 2208
rect 3744 2148 3748 2204
rect 3748 2148 3804 2204
rect 3804 2148 3808 2204
rect 3744 2144 3808 2148
rect 3824 2204 3888 2208
rect 3824 2148 3828 2204
rect 3828 2148 3884 2204
rect 3884 2148 3888 2204
rect 3824 2144 3888 2148
rect 3904 2204 3968 2208
rect 3904 2148 3908 2204
rect 3908 2148 3964 2204
rect 3964 2148 3968 2204
rect 3904 2144 3968 2148
rect 4324 1660 4388 1664
rect 4324 1604 4328 1660
rect 4328 1604 4384 1660
rect 4384 1604 4388 1660
rect 4324 1600 4388 1604
rect 4404 1660 4468 1664
rect 4404 1604 4408 1660
rect 4408 1604 4464 1660
rect 4464 1604 4468 1660
rect 4404 1600 4468 1604
rect 4484 1660 4548 1664
rect 4484 1604 4488 1660
rect 4488 1604 4544 1660
rect 4544 1604 4548 1660
rect 4484 1600 4548 1604
rect 4564 1660 4628 1664
rect 4564 1604 4568 1660
rect 4568 1604 4624 1660
rect 4624 1604 4628 1660
rect 4564 1600 4628 1604
rect 3664 1116 3728 1120
rect 3664 1060 3668 1116
rect 3668 1060 3724 1116
rect 3724 1060 3728 1116
rect 3664 1056 3728 1060
rect 3744 1116 3808 1120
rect 3744 1060 3748 1116
rect 3748 1060 3804 1116
rect 3804 1060 3808 1116
rect 3744 1056 3808 1060
rect 3824 1116 3888 1120
rect 3824 1060 3828 1116
rect 3828 1060 3884 1116
rect 3884 1060 3888 1116
rect 3824 1056 3888 1060
rect 3904 1116 3968 1120
rect 3904 1060 3908 1116
rect 3908 1060 3964 1116
rect 3964 1060 3968 1116
rect 3904 1056 3968 1060
rect 4324 572 4388 576
rect 4324 516 4328 572
rect 4328 516 4384 572
rect 4384 516 4388 572
rect 4324 512 4388 516
rect 4404 572 4468 576
rect 4404 516 4408 572
rect 4408 516 4464 572
rect 4464 516 4468 572
rect 4404 512 4468 516
rect 4484 572 4548 576
rect 4484 516 4488 572
rect 4488 516 4544 572
rect 4544 516 4548 572
rect 4484 512 4548 516
rect 4564 572 4628 576
rect 4564 516 4568 572
rect 4568 516 4624 572
rect 4624 516 4628 572
rect 4564 512 4628 516
<< metal4 >>
rect 3656 22880 3976 23440
rect 3656 22816 3664 22880
rect 3728 22816 3744 22880
rect 3808 22816 3824 22880
rect 3888 22816 3904 22880
rect 3968 22816 3976 22880
rect 3656 21792 3976 22816
rect 3656 21728 3664 21792
rect 3728 21728 3744 21792
rect 3808 21728 3824 21792
rect 3888 21728 3904 21792
rect 3968 21728 3976 21792
rect 3656 20704 3976 21728
rect 3656 20640 3664 20704
rect 3728 20640 3744 20704
rect 3808 20640 3824 20704
rect 3888 20640 3904 20704
rect 3968 20640 3976 20704
rect 3656 19616 3976 20640
rect 3656 19552 3664 19616
rect 3728 19552 3744 19616
rect 3808 19552 3824 19616
rect 3888 19552 3904 19616
rect 3968 19552 3976 19616
rect 3656 18528 3976 19552
rect 3656 18464 3664 18528
rect 3728 18464 3744 18528
rect 3808 18464 3824 18528
rect 3888 18464 3904 18528
rect 3968 18464 3976 18528
rect 3656 17440 3976 18464
rect 3656 17376 3664 17440
rect 3728 17376 3744 17440
rect 3808 17376 3824 17440
rect 3888 17376 3904 17440
rect 3968 17376 3976 17440
rect 3656 16352 3976 17376
rect 3656 16288 3664 16352
rect 3728 16288 3744 16352
rect 3808 16288 3824 16352
rect 3888 16288 3904 16352
rect 3968 16288 3976 16352
rect 3656 15264 3976 16288
rect 3656 15200 3664 15264
rect 3728 15200 3744 15264
rect 3808 15200 3824 15264
rect 3888 15200 3904 15264
rect 3968 15200 3976 15264
rect 3656 14176 3976 15200
rect 3656 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3904 14176
rect 3968 14112 3976 14176
rect 3656 13088 3976 14112
rect 3656 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3904 13088
rect 3968 13024 3976 13088
rect 3656 12000 3976 13024
rect 3656 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3904 12000
rect 3968 11936 3976 12000
rect 3656 10912 3976 11936
rect 3656 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3904 10912
rect 3968 10848 3976 10912
rect 3656 9824 3976 10848
rect 3656 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3904 9824
rect 3968 9760 3976 9824
rect 3656 8736 3976 9760
rect 3656 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3904 8736
rect 3968 8672 3976 8736
rect 3656 7648 3976 8672
rect 3656 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3904 7648
rect 3968 7584 3976 7648
rect 3656 6560 3976 7584
rect 3656 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3976 6560
rect 3656 5472 3976 6496
rect 3656 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3976 5472
rect 3656 4384 3976 5408
rect 3656 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3976 4384
rect 3656 3296 3976 4320
rect 3656 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3976 3296
rect 3656 2208 3976 3232
rect 3656 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3976 2208
rect 3656 1120 3976 2144
rect 3656 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3976 1120
rect 3656 496 3976 1056
rect 4316 23424 4636 23440
rect 4316 23360 4324 23424
rect 4388 23360 4404 23424
rect 4468 23360 4484 23424
rect 4548 23360 4564 23424
rect 4628 23360 4636 23424
rect 4316 22336 4636 23360
rect 4316 22272 4324 22336
rect 4388 22272 4404 22336
rect 4468 22272 4484 22336
rect 4548 22272 4564 22336
rect 4628 22272 4636 22336
rect 4316 21248 4636 22272
rect 4316 21184 4324 21248
rect 4388 21184 4404 21248
rect 4468 21184 4484 21248
rect 4548 21184 4564 21248
rect 4628 21184 4636 21248
rect 4316 20160 4636 21184
rect 4316 20096 4324 20160
rect 4388 20096 4404 20160
rect 4468 20096 4484 20160
rect 4548 20096 4564 20160
rect 4628 20096 4636 20160
rect 4316 19072 4636 20096
rect 4316 19008 4324 19072
rect 4388 19008 4404 19072
rect 4468 19008 4484 19072
rect 4548 19008 4564 19072
rect 4628 19008 4636 19072
rect 4316 17984 4636 19008
rect 4316 17920 4324 17984
rect 4388 17920 4404 17984
rect 4468 17920 4484 17984
rect 4548 17920 4564 17984
rect 4628 17920 4636 17984
rect 4316 16896 4636 17920
rect 4316 16832 4324 16896
rect 4388 16832 4404 16896
rect 4468 16832 4484 16896
rect 4548 16832 4564 16896
rect 4628 16832 4636 16896
rect 4316 15808 4636 16832
rect 4316 15744 4324 15808
rect 4388 15744 4404 15808
rect 4468 15744 4484 15808
rect 4548 15744 4564 15808
rect 4628 15744 4636 15808
rect 4316 14720 4636 15744
rect 4316 14656 4324 14720
rect 4388 14656 4404 14720
rect 4468 14656 4484 14720
rect 4548 14656 4564 14720
rect 4628 14656 4636 14720
rect 4316 13632 4636 14656
rect 4316 13568 4324 13632
rect 4388 13568 4404 13632
rect 4468 13568 4484 13632
rect 4548 13568 4564 13632
rect 4628 13568 4636 13632
rect 4316 12544 4636 13568
rect 4316 12480 4324 12544
rect 4388 12480 4404 12544
rect 4468 12480 4484 12544
rect 4548 12480 4564 12544
rect 4628 12480 4636 12544
rect 4316 11456 4636 12480
rect 4316 11392 4324 11456
rect 4388 11392 4404 11456
rect 4468 11392 4484 11456
rect 4548 11392 4564 11456
rect 4628 11392 4636 11456
rect 4316 10368 4636 11392
rect 4316 10304 4324 10368
rect 4388 10304 4404 10368
rect 4468 10304 4484 10368
rect 4548 10304 4564 10368
rect 4628 10304 4636 10368
rect 4316 9280 4636 10304
rect 4316 9216 4324 9280
rect 4388 9216 4404 9280
rect 4468 9216 4484 9280
rect 4548 9216 4564 9280
rect 4628 9216 4636 9280
rect 4316 8192 4636 9216
rect 4316 8128 4324 8192
rect 4388 8128 4404 8192
rect 4468 8128 4484 8192
rect 4548 8128 4564 8192
rect 4628 8128 4636 8192
rect 4316 7104 4636 8128
rect 4316 7040 4324 7104
rect 4388 7040 4404 7104
rect 4468 7040 4484 7104
rect 4548 7040 4564 7104
rect 4628 7040 4636 7104
rect 4316 6016 4636 7040
rect 4316 5952 4324 6016
rect 4388 5952 4404 6016
rect 4468 5952 4484 6016
rect 4548 5952 4564 6016
rect 4628 5952 4636 6016
rect 4316 4928 4636 5952
rect 4316 4864 4324 4928
rect 4388 4864 4404 4928
rect 4468 4864 4484 4928
rect 4548 4864 4564 4928
rect 4628 4864 4636 4928
rect 4316 3840 4636 4864
rect 4316 3776 4324 3840
rect 4388 3776 4404 3840
rect 4468 3776 4484 3840
rect 4548 3776 4564 3840
rect 4628 3776 4636 3840
rect 4316 2752 4636 3776
rect 4316 2688 4324 2752
rect 4388 2688 4404 2752
rect 4468 2688 4484 2752
rect 4548 2688 4564 2752
rect 4628 2688 4636 2752
rect 4316 1664 4636 2688
rect 4316 1600 4324 1664
rect 4388 1600 4404 1664
rect 4468 1600 4484 1664
rect 4548 1600 4564 1664
rect 4628 1600 4636 1664
rect 4316 576 4636 1600
rect 4316 512 4324 576
rect 4388 512 4404 576
rect 4468 512 4484 576
rect 4548 512 4564 576
rect 4628 512 4636 576
rect 4316 496 4636 512
use sky130_fd_sc_hd__inv_2  _0490_
timestamp 1729294469
transform 1 0 22724 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0491_
timestamp 1729294469
transform 1 0 20884 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0492_
timestamp 1729294469
transform 1 0 4048 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0493_
timestamp 1729294469
transform 1 0 2852 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0494_
timestamp 1729294469
transform -1 0 7084 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_6  _0495_
timestamp 1729294469
transform -1 0 21896 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0496_
timestamp 1729294469
transform 1 0 4324 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0497_
timestamp 1729294469
transform 1 0 4600 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0498_
timestamp 1729294469
transform 1 0 7728 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0499_
timestamp 1729294469
transform 1 0 8372 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0500_
timestamp 1729294469
transform -1 0 10672 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0501_
timestamp 1729294469
transform 1 0 11408 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0502_
timestamp 1729294469
transform -1 0 13432 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0503_
timestamp 1729294469
transform 1 0 14076 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0504_
timestamp 1729294469
transform 1 0 16008 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0505_
timestamp 1729294469
transform 1 0 17296 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0506_
timestamp 1729294469
transform 1 0 18952 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0507_
timestamp 1729294469
transform 1 0 19872 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _0508_
timestamp 1729294469
transform 1 0 22172 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0509_
timestamp 1729294469
transform 1 0 21804 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_4  _0510_
timestamp 1729294469
transform 1 0 21988 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  _0511_
timestamp 1729294469
transform -1 0 3864 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0512_
timestamp 1729294469
transform 1 0 2668 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0513_
timestamp 1729294469
transform -1 0 3128 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0514_
timestamp 1729294469
transform 1 0 3220 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0515_
timestamp 1729294469
transform 1 0 2760 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _0516_
timestamp 1729294469
transform -1 0 3220 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0517_
timestamp 1729294469
transform 1 0 2576 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0518_
timestamp 1729294469
transform 1 0 3864 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0519_
timestamp 1729294469
transform 1 0 4692 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0520_
timestamp 1729294469
transform 1 0 2668 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _0521_
timestamp 1729294469
transform 1 0 3956 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0522_
timestamp 1729294469
transform 1 0 4140 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0523_
timestamp 1729294469
transform 1 0 4508 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0524_
timestamp 1729294469
transform -1 0 9384 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0525_
timestamp 1729294469
transform -1 0 9476 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _0526_
timestamp 1729294469
transform -1 0 6164 0 1 22304
box -38 -48 2062 592
use sky130_fd_sc_hd__mux2_1  _0527_
timestamp 1729294469
transform 1 0 5980 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0528_
timestamp 1729294469
transform 1 0 5796 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__and3_2  _0529_
timestamp 1729294469
transform 1 0 3312 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  _0530_
timestamp 1729294469
transform 1 0 3404 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0531_
timestamp 1729294469
transform -1 0 6072 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0532_
timestamp 1729294469
transform -1 0 8280 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0533_
timestamp 1729294469
transform 1 0 8372 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0534_
timestamp 1729294469
transform 1 0 6256 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0535_
timestamp 1729294469
transform 1 0 8372 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _0536_
timestamp 1729294469
transform -1 0 5704 0 -1 21216
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _0537_
timestamp 1729294469
transform 1 0 3680 0 -1 22304
box -38 -48 2062 592
use sky130_fd_sc_hd__a21boi_2  _0538_
timestamp 1729294469
transform 1 0 3220 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _0539_
timestamp 1729294469
transform -1 0 4324 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0540_
timestamp 1729294469
transform 1 0 5060 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _0541_
timestamp 1729294469
transform 1 0 4508 0 -1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0542_
timestamp 1729294469
transform 1 0 7544 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0543_
timestamp 1729294469
transform 1 0 6992 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0544_
timestamp 1729294469
transform 1 0 7820 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0545_
timestamp 1729294469
transform -1 0 7728 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0546_
timestamp 1729294469
transform 1 0 7268 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0547_
timestamp 1729294469
transform 1 0 6624 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0548_
timestamp 1729294469
transform -1 0 7544 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0549_
timestamp 1729294469
transform -1 0 7544 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0550_
timestamp 1729294469
transform 1 0 8004 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0551_
timestamp 1729294469
transform 1 0 6992 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0552_
timestamp 1729294469
transform -1 0 7636 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _0553_
timestamp 1729294469
transform -1 0 8832 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0554_
timestamp 1729294469
transform 1 0 10304 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _0555_
timestamp 1729294469
transform -1 0 11500 0 1 19040
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _0556_
timestamp 1729294469
transform -1 0 8832 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0557_
timestamp 1729294469
transform 1 0 3588 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0558_
timestamp 1729294469
transform 1 0 4416 0 -1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_2  _0559_
timestamp 1729294469
transform -1 0 4876 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0560_
timestamp 1729294469
transform -1 0 6532 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0561_
timestamp 1729294469
transform 1 0 5980 0 -1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0562_
timestamp 1729294469
transform 1 0 7636 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0563_
timestamp 1729294469
transform -1 0 8648 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0564_
timestamp 1729294469
transform 1 0 8188 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0565_
timestamp 1729294469
transform -1 0 8740 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0566_
timestamp 1729294469
transform 1 0 8372 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0567_
timestamp 1729294469
transform -1 0 8188 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0568_
timestamp 1729294469
transform 1 0 8004 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0569_
timestamp 1729294469
transform 1 0 7636 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0570_
timestamp 1729294469
transform 1 0 8372 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_4  _0571_
timestamp 1729294469
transform -1 0 10304 0 -1 19040
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _0572_
timestamp 1729294469
transform -1 0 9660 0 -1 20128
box -38 -48 2062 592
use sky130_fd_sc_hd__a21boi_1  _0573_
timestamp 1729294469
transform 1 0 2944 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0574_
timestamp 1729294469
transform 1 0 4600 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0575_
timestamp 1729294469
transform 1 0 3680 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _0576_
timestamp 1729294469
transform 1 0 3772 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0577_
timestamp 1729294469
transform 1 0 5244 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0578_
timestamp 1729294469
transform 1 0 4968 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0579_
timestamp 1729294469
transform 1 0 5888 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0580_
timestamp 1729294469
transform 1 0 8372 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _0581_
timestamp 1729294469
transform -1 0 8280 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0582_
timestamp 1729294469
transform 1 0 7820 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0583_
timestamp 1729294469
transform 1 0 9200 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0584_
timestamp 1729294469
transform -1 0 9292 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0585_
timestamp 1729294469
transform 1 0 9200 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0586_
timestamp 1729294469
transform 1 0 8832 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0587_
timestamp 1729294469
transform -1 0 9568 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0588_
timestamp 1729294469
transform -1 0 8924 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0589_
timestamp 1729294469
transform 1 0 8924 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0590_
timestamp 1729294469
transform 1 0 10028 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _0591_
timestamp 1729294469
transform 1 0 9200 0 1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _0592_
timestamp 1729294469
transform -1 0 4784 0 1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__o31a_1  _0593_
timestamp 1729294469
transform -1 0 3864 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0594_
timestamp 1729294469
transform 1 0 3312 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0595_
timestamp 1729294469
transform -1 0 4232 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0596_
timestamp 1729294469
transform 1 0 4324 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0597_
timestamp 1729294469
transform 1 0 3956 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0598_
timestamp 1729294469
transform 1 0 5796 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0599_
timestamp 1729294469
transform -1 0 6348 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _0600_
timestamp 1729294469
transform 1 0 7176 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0601_
timestamp 1729294469
transform 1 0 6532 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0602_
timestamp 1729294469
transform 1 0 10580 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0603_
timestamp 1729294469
transform 1 0 9476 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0604_
timestamp 1729294469
transform 1 0 9476 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0605_
timestamp 1729294469
transform 1 0 10488 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0606_
timestamp 1729294469
transform -1 0 10488 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _0607_
timestamp 1729294469
transform 1 0 8464 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0608_
timestamp 1729294469
transform -1 0 8280 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0609_
timestamp 1729294469
transform 1 0 10120 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _0610_
timestamp 1729294469
transform 1 0 9384 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0611_
timestamp 1729294469
transform 1 0 10028 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0612_
timestamp 1729294469
transform 1 0 10396 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0613_
timestamp 1729294469
transform 1 0 10396 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0614_
timestamp 1729294469
transform -1 0 15272 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0615_
timestamp 1729294469
transform 1 0 15272 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0616_
timestamp 1729294469
transform -1 0 15732 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0617_
timestamp 1729294469
transform -1 0 15272 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0618_
timestamp 1729294469
transform 1 0 15180 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0619_
timestamp 1729294469
transform -1 0 14352 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_2  _0620_
timestamp 1729294469
transform 1 0 7268 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _0621_
timestamp 1729294469
transform -1 0 7912 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0622_
timestamp 1729294469
transform -1 0 9016 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0623_
timestamp 1729294469
transform -1 0 7820 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0624_
timestamp 1729294469
transform 1 0 10396 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0625_
timestamp 1729294469
transform 1 0 9936 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _0626_
timestamp 1729294469
transform 1 0 5336 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0627_
timestamp 1729294469
transform -1 0 12052 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0628_
timestamp 1729294469
transform -1 0 11592 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0629_
timestamp 1729294469
transform 1 0 10764 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0630_
timestamp 1729294469
transform -1 0 11776 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0631_
timestamp 1729294469
transform 1 0 11776 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0632_
timestamp 1729294469
transform -1 0 12880 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0633_
timestamp 1729294469
transform -1 0 12604 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0634_
timestamp 1729294469
transform 1 0 11684 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2ai_1  _0635_
timestamp 1729294469
transform 1 0 11224 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0636_
timestamp 1729294469
transform -1 0 13984 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_4  _0637_
timestamp 1729294469
transform 1 0 16100 0 -1 22304
box -38 -48 1418 592
use sky130_fd_sc_hd__a21oi_2  _0638_
timestamp 1729294469
transform 1 0 17848 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0639_
timestamp 1729294469
transform 1 0 17388 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0640_
timestamp 1729294469
transform 1 0 18308 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0641_
timestamp 1729294469
transform 1 0 18676 0 1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__a211o_1  _0642_
timestamp 1729294469
transform -1 0 7360 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_2  _0643_
timestamp 1729294469
transform -1 0 8280 0 -1 22304
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0644_
timestamp 1729294469
transform -1 0 13800 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0645_
timestamp 1729294469
transform -1 0 12144 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0646_
timestamp 1729294469
transform -1 0 10580 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0647_
timestamp 1729294469
transform -1 0 12696 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0648_
timestamp 1729294469
transform -1 0 14168 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0649_
timestamp 1729294469
transform 1 0 12236 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _0650_
timestamp 1729294469
transform 1 0 12972 0 -1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _0651_
timestamp 1729294469
transform -1 0 11500 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0652_
timestamp 1729294469
transform 1 0 13524 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _0653_
timestamp 1729294469
transform -1 0 13432 0 1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _0654_
timestamp 1729294469
transform -1 0 13800 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0655_
timestamp 1729294469
transform 1 0 12880 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0656_
timestamp 1729294469
transform 1 0 13064 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _0657_
timestamp 1729294469
transform 1 0 12236 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_4  _0658_
timestamp 1729294469
transform 1 0 18124 0 -1 22304
box -38 -48 1418 592
use sky130_fd_sc_hd__nor2_1  _0659_
timestamp 1729294469
transform 1 0 9200 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0660_
timestamp 1729294469
transform 1 0 8924 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0661_
timestamp 1729294469
transform 1 0 9844 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0662_
timestamp 1729294469
transform 1 0 4784 0 1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _0663_
timestamp 1729294469
transform 1 0 9384 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0664_
timestamp 1729294469
transform 1 0 9200 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _0665_
timestamp 1729294469
transform 1 0 10948 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__a21boi_1  _0666_
timestamp 1729294469
transform 1 0 11684 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0667_
timestamp 1729294469
transform 1 0 12696 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _0668_
timestamp 1729294469
transform 1 0 12144 0 -1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _0669_
timestamp 1729294469
transform -1 0 14720 0 1 21216
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0670_
timestamp 1729294469
transform -1 0 14352 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0671_
timestamp 1729294469
transform -1 0 13432 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0672_
timestamp 1729294469
transform -1 0 13524 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0673_
timestamp 1729294469
transform -1 0 14260 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0674_
timestamp 1729294469
transform 1 0 14260 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0675_
timestamp 1729294469
transform -1 0 13892 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0676_
timestamp 1729294469
transform 1 0 14168 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0677_
timestamp 1729294469
transform -1 0 5796 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _0678_
timestamp 1729294469
transform 1 0 6256 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0679_
timestamp 1729294469
transform 1 0 9660 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0680_
timestamp 1729294469
transform -1 0 11132 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0681_
timestamp 1729294469
transform 1 0 11224 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0682_
timestamp 1729294469
transform 1 0 10948 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0683_
timestamp 1729294469
transform 1 0 11960 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0684_
timestamp 1729294469
transform 1 0 11776 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _0685_
timestamp 1729294469
transform 1 0 12696 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _0686_
timestamp 1729294469
transform 1 0 12972 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0687_
timestamp 1729294469
transform 1 0 12788 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0688_
timestamp 1729294469
transform -1 0 14168 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0689_
timestamp 1729294469
transform 1 0 13524 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0690_
timestamp 1729294469
transform -1 0 13984 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0691_
timestamp 1729294469
transform 1 0 13524 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0692_
timestamp 1729294469
transform 1 0 13616 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0693_
timestamp 1729294469
transform 1 0 8372 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0694_
timestamp 1729294469
transform 1 0 6440 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0695_
timestamp 1729294469
transform 1 0 10028 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0696_
timestamp 1729294469
transform 1 0 9384 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0697_
timestamp 1729294469
transform 1 0 11316 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0698_
timestamp 1729294469
transform -1 0 12972 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0699_
timestamp 1729294469
transform 1 0 12512 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0700_
timestamp 1729294469
transform 1 0 12880 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0701_
timestamp 1729294469
transform 1 0 13892 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0702_
timestamp 1729294469
transform -1 0 14720 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0703_
timestamp 1729294469
transform 1 0 13524 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0704_
timestamp 1729294469
transform 1 0 14904 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0705_
timestamp 1729294469
transform 1 0 3128 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0706_
timestamp 1729294469
transform 1 0 4416 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0707_
timestamp 1729294469
transform -1 0 6164 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0708_
timestamp 1729294469
transform 1 0 5612 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0709_
timestamp 1729294469
transform 1 0 6992 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _0710_
timestamp 1729294469
transform -1 0 8280 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0711_
timestamp 1729294469
transform 1 0 9752 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0712_
timestamp 1729294469
transform 1 0 9108 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0713_
timestamp 1729294469
transform 1 0 10212 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_2  _0714_
timestamp 1729294469
transform 1 0 10396 0 1 17952
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0715_
timestamp 1729294469
transform 1 0 12420 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1729294469
transform 1 0 16744 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0717_
timestamp 1729294469
transform 1 0 11776 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0718_
timestamp 1729294469
transform 1 0 13064 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0719_
timestamp 1729294469
transform -1 0 14076 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0720_
timestamp 1729294469
transform -1 0 13892 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0721_
timestamp 1729294469
transform 1 0 15548 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0722_
timestamp 1729294469
transform -1 0 15548 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0723_
timestamp 1729294469
transform -1 0 16008 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0724_
timestamp 1729294469
transform 1 0 4784 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0725_
timestamp 1729294469
transform 1 0 4140 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0726_
timestamp 1729294469
transform 1 0 4692 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0727_
timestamp 1729294469
transform -1 0 4508 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0728_
timestamp 1729294469
transform 1 0 5152 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0729_
timestamp 1729294469
transform 1 0 4784 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0730_
timestamp 1729294469
transform 1 0 5796 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0731_
timestamp 1729294469
transform -1 0 7728 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0732_
timestamp 1729294469
transform 1 0 15732 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0733_
timestamp 1729294469
transform 1 0 14444 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0734_
timestamp 1729294469
transform 1 0 15088 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_2  _0735_
timestamp 1729294469
transform 1 0 10948 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0736_
timestamp 1729294469
transform 1 0 15640 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0737_
timestamp 1729294469
transform 1 0 15088 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0738_
timestamp 1729294469
transform 1 0 15364 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1729294469
transform 1 0 16468 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0740_
timestamp 1729294469
transform 1 0 16560 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0741_
timestamp 1729294469
transform -1 0 16560 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0742_
timestamp 1729294469
transform -1 0 16744 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0743_
timestamp 1729294469
transform 1 0 14720 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0744_
timestamp 1729294469
transform 1 0 14720 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0745_
timestamp 1729294469
transform -1 0 15640 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0746_
timestamp 1729294469
transform 1 0 16008 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0747_
timestamp 1729294469
transform 1 0 15732 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0748_
timestamp 1729294469
transform -1 0 16652 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0749_
timestamp 1729294469
transform -1 0 6256 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0750_
timestamp 1729294469
transform 1 0 16468 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0751_
timestamp 1729294469
transform 1 0 15824 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0752_
timestamp 1729294469
transform 1 0 16928 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0753_
timestamp 1729294469
transform 1 0 16284 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0754_
timestamp 1729294469
transform -1 0 16560 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0755_
timestamp 1729294469
transform -1 0 17480 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0756_
timestamp 1729294469
transform 1 0 17204 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0757_
timestamp 1729294469
transform 1 0 17664 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _0758_
timestamp 1729294469
transform -1 0 13248 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _0759_
timestamp 1729294469
transform -1 0 16008 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _0760_
timestamp 1729294469
transform 1 0 14168 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0761_
timestamp 1729294469
transform 1 0 16008 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0762_
timestamp 1729294469
transform -1 0 16836 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0763_
timestamp 1729294469
transform 1 0 17020 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0764_
timestamp 1729294469
transform 1 0 18216 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0765_
timestamp 1729294469
transform -1 0 18124 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0766_
timestamp 1729294469
transform 1 0 18676 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _0767_
timestamp 1729294469
transform 1 0 17940 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0768_
timestamp 1729294469
transform 1 0 16560 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0769_
timestamp 1729294469
transform -1 0 17112 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0770_
timestamp 1729294469
transform 1 0 17204 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0771_
timestamp 1729294469
transform 1 0 17664 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1729294469
transform 1 0 17664 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0773_
timestamp 1729294469
transform 1 0 17204 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0774_
timestamp 1729294469
transform 1 0 17296 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0775_
timestamp 1729294469
transform -1 0 17940 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0776_
timestamp 1729294469
transform -1 0 18308 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0777_
timestamp 1729294469
transform 1 0 18124 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0778_
timestamp 1729294469
transform 1 0 18676 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0779_
timestamp 1729294469
transform 1 0 18676 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0780_
timestamp 1729294469
transform -1 0 21528 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0781_
timestamp 1729294469
transform -1 0 20700 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0782_
timestamp 1729294469
transform 1 0 19872 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0783_
timestamp 1729294469
transform -1 0 21988 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0784_
timestamp 1729294469
transform 1 0 20424 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0785_
timestamp 1729294469
transform 1 0 20332 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0786_
timestamp 1729294469
transform 1 0 20884 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0787_
timestamp 1729294469
transform -1 0 18492 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _0788_
timestamp 1729294469
transform 1 0 19504 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0789_
timestamp 1729294469
transform -1 0 19780 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0790_
timestamp 1729294469
transform -1 0 19688 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__o311ai_2  _0791_
timestamp 1729294469
transform 1 0 17020 0 -1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0792_
timestamp 1729294469
transform 1 0 18308 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0793_
timestamp 1729294469
transform -1 0 18400 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0794_
timestamp 1729294469
transform -1 0 19228 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0795_
timestamp 1729294469
transform 1 0 18860 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0796_
timestamp 1729294469
transform -1 0 20148 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0797_
timestamp 1729294469
transform 1 0 19228 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0798_
timestamp 1729294469
transform -1 0 22816 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0799_
timestamp 1729294469
transform -1 0 22080 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _0800_
timestamp 1729294469
transform -1 0 21528 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _0801_
timestamp 1729294469
transform 1 0 21896 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0802_
timestamp 1729294469
transform -1 0 22448 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0803_
timestamp 1729294469
transform -1 0 20884 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0804_
timestamp 1729294469
transform -1 0 21804 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0805_
timestamp 1729294469
transform -1 0 21344 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0806_
timestamp 1729294469
transform -1 0 20424 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0807_
timestamp 1729294469
transform 1 0 21252 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _0808_
timestamp 1729294469
transform 1 0 21252 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0809_
timestamp 1729294469
transform 1 0 20608 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0810_
timestamp 1729294469
transform 1 0 20332 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0811_
timestamp 1729294469
transform -1 0 21712 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0812_
timestamp 1729294469
transform 1 0 19872 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0813_
timestamp 1729294469
transform 1 0 21252 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0814_
timestamp 1729294469
transform 1 0 21436 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0815_
timestamp 1729294469
transform 1 0 22172 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0816_
timestamp 1729294469
transform 1 0 20424 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0817_
timestamp 1729294469
transform 1 0 21252 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0818_
timestamp 1729294469
transform 1 0 21712 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0819_
timestamp 1729294469
transform 1 0 21528 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0820_
timestamp 1729294469
transform 1 0 20976 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0821_
timestamp 1729294469
transform 1 0 21344 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0822_
timestamp 1729294469
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0823_
timestamp 1729294469
transform -1 0 21160 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0824_
timestamp 1729294469
transform 1 0 20148 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0825_
timestamp 1729294469
transform 1 0 19412 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0826_
timestamp 1729294469
transform 1 0 19780 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0827_
timestamp 1729294469
transform 1 0 19320 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0828_
timestamp 1729294469
transform -1 0 19320 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0829_
timestamp 1729294469
transform -1 0 18676 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0830_
timestamp 1729294469
transform 1 0 17204 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0831_
timestamp 1729294469
transform 1 0 17480 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0832_
timestamp 1729294469
transform -1 0 18032 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0833_
timestamp 1729294469
transform 1 0 18676 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0834_
timestamp 1729294469
transform 1 0 16468 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0835_
timestamp 1729294469
transform 1 0 16652 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0836_
timestamp 1729294469
transform -1 0 17480 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0837_
timestamp 1729294469
transform 1 0 17296 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0838_
timestamp 1729294469
transform 1 0 15364 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0839_
timestamp 1729294469
transform 1 0 16100 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _0840_
timestamp 1729294469
transform 1 0 12880 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0841_
timestamp 1729294469
transform 1 0 15548 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0842_
timestamp 1729294469
transform -1 0 15916 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0843_
timestamp 1729294469
transform 1 0 13524 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0844_
timestamp 1729294469
transform -1 0 14812 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0845_
timestamp 1729294469
transform -1 0 14628 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0846_
timestamp 1729294469
transform -1 0 13800 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0847_
timestamp 1729294469
transform 1 0 13524 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _0848_
timestamp 1729294469
transform 1 0 11132 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0849_
timestamp 1729294469
transform 1 0 12328 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0850_
timestamp 1729294469
transform 1 0 12696 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0851_
timestamp 1729294469
transform -1 0 11592 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0852_
timestamp 1729294469
transform 1 0 10948 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0853_
timestamp 1729294469
transform 1 0 10672 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0854_
timestamp 1729294469
transform 1 0 11592 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0855_
timestamp 1729294469
transform 1 0 10488 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0856_
timestamp 1729294469
transform 1 0 8372 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0857_
timestamp 1729294469
transform 1 0 9384 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0858_
timestamp 1729294469
transform 1 0 7360 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0859_
timestamp 1729294469
transform -1 0 8832 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0860_
timestamp 1729294469
transform 1 0 7912 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0861_
timestamp 1729294469
transform 1 0 6348 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0862_
timestamp 1729294469
transform 1 0 6900 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0863_
timestamp 1729294469
transform 1 0 5612 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0864_
timestamp 1729294469
transform 1 0 5796 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0865_
timestamp 1729294469
transform -1 0 6624 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0866_
timestamp 1729294469
transform 1 0 4784 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0867_
timestamp 1729294469
transform 1 0 4600 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0868_
timestamp 1729294469
transform 1 0 5244 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0869_
timestamp 1729294469
transform 1 0 3128 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0870_
timestamp 1729294469
transform 1 0 3772 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0871_
timestamp 1729294469
transform -1 0 5796 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0872_
timestamp 1729294469
transform -1 0 3220 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0873_
timestamp 1729294469
transform -1 0 4508 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0874_
timestamp 1729294469
transform 1 0 3312 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0875_
timestamp 1729294469
transform -1 0 3312 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0876_
timestamp 1729294469
transform 1 0 3680 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _0877_
timestamp 1729294469
transform 1 0 4600 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0878_
timestamp 1729294469
transform 1 0 5888 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0879_
timestamp 1729294469
transform 1 0 7820 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0880_
timestamp 1729294469
transform 1 0 11592 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0881_
timestamp 1729294469
transform 1 0 13984 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0882_
timestamp 1729294469
transform 1 0 16744 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0883_
timestamp 1729294469
transform 1 0 17940 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0884_
timestamp 1729294469
transform 1 0 20148 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _0885_
timestamp 1729294469
transform -1 0 22540 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0886_
timestamp 1729294469
transform -1 0 22908 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _0887_
timestamp 1729294469
transform 1 0 21436 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0888_
timestamp 1729294469
transform 1 0 21620 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0889_
timestamp 1729294469
transform -1 0 2392 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0890_
timestamp 1729294469
transform -1 0 5152 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0891_
timestamp 1729294469
transform -1 0 4968 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0892_
timestamp 1729294469
transform 1 0 3404 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0893_
timestamp 1729294469
transform 1 0 3312 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0894_
timestamp 1729294469
transform 1 0 3220 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0895_
timestamp 1729294469
transform -1 0 3128 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0896_
timestamp 1729294469
transform 1 0 2208 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0897_
timestamp 1729294469
transform -1 0 2944 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0898_
timestamp 1729294469
transform -1 0 2576 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0899_
timestamp 1729294469
transform -1 0 3680 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0900_
timestamp 1729294469
transform 1 0 2944 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0901_
timestamp 1729294469
transform 1 0 2576 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0902_
timestamp 1729294469
transform 1 0 3772 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0903_
timestamp 1729294469
transform 1 0 4692 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0904_
timestamp 1729294469
transform 1 0 4232 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0905_
timestamp 1729294469
transform -1 0 6256 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0906_
timestamp 1729294469
transform 1 0 5244 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0907_
timestamp 1729294469
transform -1 0 5980 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0908_
timestamp 1729294469
transform -1 0 6992 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0909_
timestamp 1729294469
transform 1 0 6900 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0910_
timestamp 1729294469
transform -1 0 6900 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0911_
timestamp 1729294469
transform 1 0 6992 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0912_
timestamp 1729294469
transform 1 0 7452 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0913_
timestamp 1729294469
transform 1 0 7636 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0914_
timestamp 1729294469
transform 1 0 9108 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0915_
timestamp 1729294469
transform -1 0 9476 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0916_
timestamp 1729294469
transform 1 0 8556 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0917_
timestamp 1729294469
transform -1 0 10672 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0918_
timestamp 1729294469
transform -1 0 10672 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0919_
timestamp 1729294469
transform -1 0 10764 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0920_
timestamp 1729294469
transform 1 0 10948 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0921_
timestamp 1729294469
transform 1 0 10948 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0922_
timestamp 1729294469
transform 1 0 11592 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0923_
timestamp 1729294469
transform -1 0 13248 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0924_
timestamp 1729294469
transform -1 0 13432 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0925_
timestamp 1729294469
transform 1 0 12512 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0926_
timestamp 1729294469
transform 1 0 13616 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0927_
timestamp 1729294469
transform 1 0 14076 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0928_
timestamp 1729294469
transform -1 0 14076 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0929_
timestamp 1729294469
transform 1 0 14076 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0930_
timestamp 1729294469
transform 1 0 14720 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0931_
timestamp 1729294469
transform 1 0 14812 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0932_
timestamp 1729294469
transform 1 0 16008 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0933_
timestamp 1729294469
transform 1 0 15548 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0934_
timestamp 1729294469
transform 1 0 16008 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0935_
timestamp 1729294469
transform -1 0 17112 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0936_
timestamp 1729294469
transform 1 0 16100 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0937_
timestamp 1729294469
transform 1 0 15088 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0938_
timestamp 1729294469
transform 1 0 16376 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0939_
timestamp 1729294469
transform 1 0 15548 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0940_
timestamp 1729294469
transform 1 0 17020 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0941_
timestamp 1729294469
transform 1 0 18308 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0942_
timestamp 1729294469
transform 1 0 18676 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0943_
timestamp 1729294469
transform -1 0 19596 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0944_
timestamp 1729294469
transform 1 0 18216 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0945_
timestamp 1729294469
transform -1 0 18584 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0946_
timestamp 1729294469
transform -1 0 19320 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0947_
timestamp 1729294469
transform 1 0 19228 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0948_
timestamp 1729294469
transform -1 0 20148 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0949_
timestamp 1729294469
transform 1 0 19504 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0950_
timestamp 1729294469
transform 1 0 19412 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0951_
timestamp 1729294469
transform 1 0 19688 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0952_
timestamp 1729294469
transform 1 0 20240 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0953_
timestamp 1729294469
transform 1 0 20792 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0954_
timestamp 1729294469
transform -1 0 21068 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0955_
timestamp 1729294469
transform 1 0 21252 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0956_
timestamp 1729294469
transform 1 0 20424 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0957_
timestamp 1729294469
transform 1 0 20884 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0958_
timestamp 1729294469
transform -1 0 21896 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0959_
timestamp 1729294469
transform -1 0 22356 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0960_
timestamp 1729294469
transform 1 0 22356 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0961_
timestamp 1729294469
transform -1 0 21896 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0962_
timestamp 1729294469
transform -1 0 22172 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0963_
timestamp 1729294469
transform 1 0 21896 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0964_
timestamp 1729294469
transform 1 0 20976 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0965_
timestamp 1729294469
transform 1 0 22172 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0966_
timestamp 1729294469
transform -1 0 20976 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0967_
timestamp 1729294469
transform 1 0 20792 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0968_
timestamp 1729294469
transform 1 0 20700 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0969_
timestamp 1729294469
transform 1 0 19964 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0970_
timestamp 1729294469
transform 1 0 20056 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0971_
timestamp 1729294469
transform -1 0 20240 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0972_
timestamp 1729294469
transform -1 0 19412 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0973_
timestamp 1729294469
transform -1 0 20148 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0974_
timestamp 1729294469
transform -1 0 19780 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0975_
timestamp 1729294469
transform -1 0 19320 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0976_
timestamp 1729294469
transform -1 0 19688 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0977_
timestamp 1729294469
transform 1 0 18308 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0978_
timestamp 1729294469
transform -1 0 19228 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0979_
timestamp 1729294469
transform -1 0 22172 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0980_
timestamp 1729294469
transform 1 0 21620 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _0981_
timestamp 1729294469
transform -1 0 4692 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0982_
timestamp 1729294469
transform -1 0 4416 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0983_
timestamp 1729294469
transform 1 0 3220 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0984_
timestamp 1729294469
transform 1 0 3956 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0985_
timestamp 1729294469
transform 1 0 5336 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0986_
timestamp 1729294469
transform 1 0 6532 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0987_
timestamp 1729294469
transform 1 0 7728 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0988_
timestamp 1729294469
transform 1 0 9384 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0989_
timestamp 1729294469
transform 1 0 9568 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0990_
timestamp 1729294469
transform 1 0 11040 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0991_
timestamp 1729294469
transform -1 0 14996 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0992_
timestamp 1729294469
transform -1 0 14168 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0993_
timestamp 1729294469
transform 1 0 13524 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0994_
timestamp 1729294469
transform 1 0 14536 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0995_
timestamp 1729294469
transform 1 0 15272 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0996_
timestamp 1729294469
transform 1 0 16744 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0997_
timestamp 1729294469
transform 1 0 18216 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0998_
timestamp 1729294469
transform 1 0 18676 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _0999_
timestamp 1729294469
transform 1 0 18860 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1000_
timestamp 1729294469
transform 1 0 20424 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1001_
timestamp 1729294469
transform 1 0 21620 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1002_
timestamp 1729294469
transform -1 0 22724 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1003_
timestamp 1729294469
transform 1 0 1656 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1004_
timestamp 1729294469
transform 1 0 4048 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1005_
timestamp 1729294469
transform 1 0 3220 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1006_
timestamp 1729294469
transform 1 0 2392 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1007_
timestamp 1729294469
transform 1 0 1656 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1008_
timestamp 1729294469
transform 1 0 3220 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1009_
timestamp 1729294469
transform -1 0 5704 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1010_
timestamp 1729294469
transform 1 0 5428 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1011_
timestamp 1729294469
transform 1 0 6072 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1012_
timestamp 1729294469
transform -1 0 9016 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1013_
timestamp 1729294469
transform 1 0 8648 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1014_
timestamp 1729294469
transform 1 0 9476 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1015_
timestamp 1729294469
transform -1 0 12420 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1016_
timestamp 1729294469
transform 1 0 12788 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1017_
timestamp 1729294469
transform 1 0 13524 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1018_
timestamp 1729294469
transform -1 0 16560 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1019_
timestamp 1729294469
transform 1 0 16100 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1020_
timestamp 1729294469
transform 1 0 15732 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1021_
timestamp 1729294469
transform -1 0 17848 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1022_
timestamp 1729294469
transform -1 0 19596 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1023_
timestamp 1729294469
transform -1 0 18584 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1024_
timestamp 1729294469
transform -1 0 20792 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1025_
timestamp 1729294469
transform -1 0 21620 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1026_
timestamp 1729294469
transform -1 0 23092 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1027_
timestamp 1729294469
transform 1 0 21344 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1028_
timestamp 1729294469
transform 1 0 21252 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1029_
timestamp 1729294469
transform 1 0 21436 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1030_
timestamp 1729294469
transform 1 0 21436 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1031_
timestamp 1729294469
transform 1 0 19688 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1032_
timestamp 1729294469
transform 1 0 18584 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1033_
timestamp 1729294469
transform 1 0 18308 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1034_
timestamp 1729294469
transform 1 0 18676 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1035_
timestamp 1729294469
transform 1 0 21436 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  fanout11
timestamp 1729294469
transform -1 0 8280 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout12
timestamp 1729294469
transform -1 0 21068 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout13
timestamp 1729294469
transform -1 0 22448 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout14
timestamp 1729294469
transform 1 0 21896 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout15
timestamp 1729294469
transform -1 0 20608 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout16
timestamp 1729294469
transform -1 0 21160 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout17
timestamp 1729294469
transform -1 0 16744 0 1 22304
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_2  fanout18
timestamp 1729294469
transform -1 0 5152 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout19
timestamp 1729294469
transform -1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout20
timestamp 1729294469
transform -1 0 3128 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout21
timestamp 1729294469
transform 1 0 19320 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout22
timestamp 1729294469
transform -1 0 22724 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout23
timestamp 1729294469
transform -1 0 6532 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout24
timestamp 1729294469
transform 1 0 9752 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout25
timestamp 1729294469
transform -1 0 11868 0 -1 4896
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout26
timestamp 1729294469
transform 1 0 20424 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout27
timestamp 1729294469
transform -1 0 21988 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout28
timestamp 1729294469
transform -1 0 23092 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout29
timestamp 1729294469
transform -1 0 22540 0 1 7072
box -38 -48 958 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 1729294469
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1729294469
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 1729294469
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1729294469
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1729294469
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 1729294469
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1729294469
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1729294469
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1729294469
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1729294469
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1729294469
transform 1 0 9476 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1729294469
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1729294469
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1729294469
transform 1 0 12052 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1729294469
transform 1 0 13156 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1729294469
transform 1 0 13524 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1729294469
transform 1 0 14628 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1729294469
transform 1 0 15732 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1729294469
transform 1 0 16100 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1729294469
transform 1 0 17204 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1729294469
transform 1 0 18308 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1729294469
transform 1 0 18676 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1729294469
transform 1 0 19780 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1729294469
transform 1 0 20884 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1729294469
transform 1 0 21252 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_237
timestamp 1729294469
transform 1 0 22356 0 1 544
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1729294469
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1729294469
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1729294469
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1729294469
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1729294469
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1729294469
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1729294469
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1729294469
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1729294469
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1729294469
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1729294469
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1729294469
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1729294469
transform 1 0 10948 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1729294469
transform 1 0 12052 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1729294469
transform 1 0 13156 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1729294469
transform 1 0 14260 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1729294469
transform 1 0 15364 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1729294469
transform 1 0 15916 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1729294469
transform 1 0 16100 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1729294469
transform 1 0 17204 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1729294469
transform 1 0 18308 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1729294469
transform 1 0 19412 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1729294469
transform 1 0 20516 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1729294469
transform 1 0 21068 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1729294469
transform 1 0 21252 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_237
timestamp 1729294469
transform 1 0 22356 0 -1 1632
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1729294469
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1729294469
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1729294469
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1729294469
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1729294469
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1729294469
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1729294469
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1729294469
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1729294469
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1729294469
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1729294469
transform 1 0 9476 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1729294469
transform 1 0 10580 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1729294469
transform 1 0 11684 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1729294469
transform 1 0 12788 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1729294469
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1729294469
transform 1 0 13524 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1729294469
transform 1 0 14628 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1729294469
transform 1 0 15732 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1729294469
transform 1 0 16836 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1729294469
transform 1 0 17940 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1729294469
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1729294469
transform 1 0 18676 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1729294469
transform 1 0 19780 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1729294469
transform 1 0 20884 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1729294469
transform 1 0 21988 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1729294469
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1729294469
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1729294469
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1729294469
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1729294469
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1729294469
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1729294469
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1729294469
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1729294469
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1729294469
transform 1 0 9108 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1729294469
transform 1 0 10212 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1729294469
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1729294469
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1729294469
transform 1 0 12052 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1729294469
transform 1 0 13156 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1729294469
transform 1 0 14260 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1729294469
transform 1 0 15364 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1729294469
transform 1 0 15916 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1729294469
transform 1 0 16100 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1729294469
transform 1 0 17204 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1729294469
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1729294469
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1729294469
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1729294469
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1729294469
transform 1 0 21252 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_237
timestamp 1729294469
transform 1 0 22356 0 -1 2720
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1729294469
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1729294469
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1729294469
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_29
timestamp 1729294469
transform 1 0 3220 0 1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_37
timestamp 1729294469
transform 1 0 3956 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_49
timestamp 1729294469
transform 1 0 5060 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_61
timestamp 1729294469
transform 1 0 6164 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_73
timestamp 1729294469
transform 1 0 7268 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_81
timestamp 1729294469
transform 1 0 8004 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1729294469
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1729294469
transform 1 0 9476 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1729294469
transform 1 0 10580 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1729294469
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1729294469
transform 1 0 12788 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1729294469
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1729294469
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1729294469
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1729294469
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1729294469
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1729294469
transform 1 0 17940 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1729294469
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1729294469
transform 1 0 18676 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1729294469
transform 1 0 19780 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1729294469
transform 1 0 20884 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1729294469
transform 1 0 21988 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1729294469
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_15
timestamp 1729294469
transform 1 0 1932 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_23
timestamp 1729294469
transform 1 0 2668 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_50
timestamp 1729294469
transform 1 0 5152 0 -1 3808
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1729294469
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1729294469
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1729294469
transform 1 0 8004 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1729294469
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1729294469
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1729294469
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1729294469
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1729294469
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1729294469
transform 1 0 13156 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1729294469
transform 1 0 14260 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1729294469
transform 1 0 15364 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1729294469
transform 1 0 15916 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1729294469
transform 1 0 16100 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1729294469
transform 1 0 17204 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1729294469
transform 1 0 18308 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1729294469
transform 1 0 19412 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1729294469
transform 1 0 20516 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1729294469
transform 1 0 21068 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1729294469
transform 1 0 21252 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_237
timestamp 1729294469
transform 1 0 22356 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_3
timestamp 1729294469
transform 1 0 828 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_11
timestamp 1729294469
transform 1 0 1564 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_36
timestamp 1729294469
transform 1 0 3864 0 1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_57
timestamp 1729294469
transform 1 0 5796 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_69
timestamp 1729294469
transform 1 0 6900 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_81
timestamp 1729294469
transform 1 0 8004 0 1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1729294469
transform 1 0 8372 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_97
timestamp 1729294469
transform 1 0 9476 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_110
timestamp 1729294469
transform 1 0 10672 0 1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_118
timestamp 1729294469
transform 1 0 11408 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_130
timestamp 1729294469
transform 1 0 12512 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_138
timestamp 1729294469
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1729294469
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1729294469
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1729294469
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1729294469
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1729294469
transform 1 0 17940 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1729294469
transform 1 0 18492 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1729294469
transform 1 0 18676 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1729294469
transform 1 0 19780 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1729294469
transform 1 0 20884 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_233
timestamp 1729294469
transform 1 0 21988 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_241
timestamp 1729294469
transform 1 0 22724 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_3
timestamp 1729294469
transform 1 0 828 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_11
timestamp 1729294469
transform 1 0 1564 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_48
timestamp 1729294469
transform 1 0 4968 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_57
timestamp 1729294469
transform 1 0 5796 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_70
timestamp 1729294469
transform 1 0 6992 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_78
timestamp 1729294469
transform 1 0 7728 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_84
timestamp 1729294469
transform 1 0 8280 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1729294469
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_123
timestamp 1729294469
transform 1 0 11868 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_131
timestamp 1729294469
transform 1 0 12604 0 -1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1729294469
transform 1 0 14260 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1729294469
transform 1 0 15364 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1729294469
transform 1 0 15916 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1729294469
transform 1 0 16100 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1729294469
transform 1 0 17204 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1729294469
transform 1 0 18308 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_205
timestamp 1729294469
transform 1 0 19412 0 -1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1729294469
transform 1 0 21252 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_237
timestamp 1729294469
transform 1 0 22356 0 -1 4896
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1729294469
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_15
timestamp 1729294469
transform 1 0 1932 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_29
timestamp 1729294469
transform 1 0 3220 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_35
timestamp 1729294469
transform 1 0 3772 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_47
timestamp 1729294469
transform 1 0 4876 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_69
timestamp 1729294469
transform 1 0 6900 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_85
timestamp 1729294469
transform 1 0 8372 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_129
timestamp 1729294469
transform 1 0 12420 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_157
timestamp 1729294469
transform 1 0 14996 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_174
timestamp 1729294469
transform 1 0 16560 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_186
timestamp 1729294469
transform 1 0 17664 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_194
timestamp 1729294469
transform 1 0 18400 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_197
timestamp 1729294469
transform 1 0 18676 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_205
timestamp 1729294469
transform 1 0 19412 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_222
timestamp 1729294469
transform 1 0 20976 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_228
timestamp 1729294469
transform 1 0 21528 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1729294469
transform 1 0 21988 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1729294469
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1729294469
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1729294469
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1729294469
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_57
timestamp 1729294469
transform 1 0 5796 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_92
timestamp 1729294469
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_96
timestamp 1729294469
transform 1 0 9384 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_110
timestamp 1729294469
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_127
timestamp 1729294469
transform 1 0 12236 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_138
timestamp 1729294469
transform 1 0 13248 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_153
timestamp 1729294469
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_162
timestamp 1729294469
transform 1 0 15456 0 -1 5984
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1729294469
transform 1 0 16100 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1729294469
transform 1 0 17204 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_193
timestamp 1729294469
transform 1 0 18308 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_218
timestamp 1729294469
transform 1 0 20608 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_240
timestamp 1729294469
transform 1 0 22632 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_244
timestamp 1729294469
transform 1 0 23000 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1729294469
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1729294469
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1729294469
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_29
timestamp 1729294469
transform 1 0 3220 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_37
timestamp 1729294469
transform 1 0 3956 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_47
timestamp 1729294469
transform 1 0 4876 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_53
timestamp 1729294469
transform 1 0 5428 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_80
timestamp 1729294469
transform 1 0 7912 0 1 5984
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1729294469
transform 1 0 8372 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1729294469
transform 1 0 9476 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1729294469
transform 1 0 10580 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1729294469
transform 1 0 11684 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1729294469
transform 1 0 12788 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1729294469
transform 1 0 13340 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_141
timestamp 1729294469
transform 1 0 13524 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_159
timestamp 1729294469
transform 1 0 15180 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_167
timestamp 1729294469
transform 1 0 15916 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_173
timestamp 1729294469
transform 1 0 16468 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_185
timestamp 1729294469
transform 1 0 17572 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_193
timestamp 1729294469
transform 1 0 18308 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_214
timestamp 1729294469
transform 1 0 20240 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_243
timestamp 1729294469
transform 1 0 22908 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1729294469
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_15
timestamp 1729294469
transform 1 0 1932 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_34
timestamp 1729294469
transform 1 0 3680 0 -1 7072
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1729294469
transform 1 0 5796 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1729294469
transform 1 0 6900 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1729294469
transform 1 0 8004 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_93
timestamp 1729294469
transform 1 0 9108 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_103
timestamp 1729294469
transform 1 0 10028 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1729294469
transform 1 0 10764 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_126
timestamp 1729294469
transform 1 0 12144 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_138
timestamp 1729294469
transform 1 0 13248 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_150
timestamp 1729294469
transform 1 0 14352 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_162
timestamp 1729294469
transform 1 0 15456 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_185
timestamp 1729294469
transform 1 0 17572 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_209
timestamp 1729294469
transform 1 0 19780 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1729294469
transform 1 0 21068 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_225
timestamp 1729294469
transform 1 0 21252 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_243
timestamp 1729294469
transform 1 0 22908 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_3
timestamp 1729294469
transform 1 0 828 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_11
timestamp 1729294469
transform 1 0 1564 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_50
timestamp 1729294469
transform 1 0 5152 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_62
timestamp 1729294469
transform 1 0 6256 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_68
timestamp 1729294469
transform 1 0 6808 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_76
timestamp 1729294469
transform 1 0 7544 0 1 7072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_90
timestamp 1729294469
transform 1 0 8832 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_102
timestamp 1729294469
transform 1 0 9936 0 1 7072
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_115
timestamp 1729294469
transform 1 0 11132 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_127
timestamp 1729294469
transform 1 0 12236 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_131
timestamp 1729294469
transform 1 0 12604 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1729294469
transform 1 0 13340 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_155
timestamp 1729294469
transform 1 0 14812 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_167
timestamp 1729294469
transform 1 0 15916 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_171
timestamp 1729294469
transform 1 0 16284 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_183
timestamp 1729294469
transform 1 0 17388 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_191
timestamp 1729294469
transform 1 0 18124 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_197
timestamp 1729294469
transform 1 0 18676 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_213
timestamp 1729294469
transform 1 0 20148 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_239
timestamp 1729294469
transform 1 0 22540 0 1 7072
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1729294469
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_15
timestamp 1729294469
transform 1 0 1932 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_32
timestamp 1729294469
transform 1 0 3496 0 -1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_42
timestamp 1729294469
transform 1 0 4416 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_54
timestamp 1729294469
transform 1 0 5520 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_57
timestamp 1729294469
transform 1 0 5796 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_70
timestamp 1729294469
transform 1 0 6992 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_78
timestamp 1729294469
transform 1 0 7728 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_92
timestamp 1729294469
transform 1 0 9016 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_104
timestamp 1729294469
transform 1 0 10120 0 -1 8160
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_123
timestamp 1729294469
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_135
timestamp 1729294469
transform 1 0 12972 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_144
timestamp 1729294469
transform 1 0 13800 0 -1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_152
timestamp 1729294469
transform 1 0 14536 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_164
timestamp 1729294469
transform 1 0 15640 0 -1 8160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_180
timestamp 1729294469
transform 1 0 17112 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_192
timestamp 1729294469
transform 1 0 18216 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_196
timestamp 1729294469
transform 1 0 18584 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_213
timestamp 1729294469
transform 1 0 20148 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_221
timestamp 1729294469
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_237
timestamp 1729294469
transform 1 0 22356 0 -1 8160
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1729294469
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1729294469
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1729294469
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_29
timestamp 1729294469
transform 1 0 3220 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_33
timestamp 1729294469
transform 1 0 3588 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_39
timestamp 1729294469
transform 1 0 4140 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_43
timestamp 1729294469
transform 1 0 4508 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_49
timestamp 1729294469
transform 1 0 5060 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_66
timestamp 1729294469
transform 1 0 6624 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1729294469
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_91
timestamp 1729294469
transform 1 0 8924 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_103
timestamp 1729294469
transform 1 0 10028 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_121
timestamp 1729294469
transform 1 0 11684 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_127
timestamp 1729294469
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_131
timestamp 1729294469
transform 1 0 12604 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_153
timestamp 1729294469
transform 1 0 14628 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_157
timestamp 1729294469
transform 1 0 14996 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_181
timestamp 1729294469
transform 1 0 17204 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_193
timestamp 1729294469
transform 1 0 18308 0 1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1729294469
transform 1 0 18676 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_209
timestamp 1729294469
transform 1 0 19780 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_221
timestamp 1729294469
transform 1 0 20884 0 1 8160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_232
timestamp 1729294469
transform 1 0 21896 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_244
timestamp 1729294469
transform 1 0 23000 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1729294469
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1729294469
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_42
timestamp 1729294469
transform 1 0 4416 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_52
timestamp 1729294469
transform 1 0 5336 0 -1 9248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1729294469
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_69
timestamp 1729294469
transform 1 0 6900 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_77
timestamp 1729294469
transform 1 0 7636 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_94
timestamp 1729294469
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_113
timestamp 1729294469
transform 1 0 10948 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_117
timestamp 1729294469
transform 1 0 11316 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1729294469
transform 1 0 12052 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_137
timestamp 1729294469
transform 1 0 13156 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_145
timestamp 1729294469
transform 1 0 13892 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_154
timestamp 1729294469
transform 1 0 14720 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_162
timestamp 1729294469
transform 1 0 15456 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_169
timestamp 1729294469
transform 1 0 16100 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_188
timestamp 1729294469
transform 1 0 17848 0 -1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_207
timestamp 1729294469
transform 1 0 19596 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_219
timestamp 1729294469
transform 1 0 20700 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1729294469
transform 1 0 21068 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_241
timestamp 1729294469
transform 1 0 22724 0 -1 9248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1729294469
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1729294469
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1729294469
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1729294469
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_41
timestamp 1729294469
transform 1 0 4324 0 1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_58
timestamp 1729294469
transform 1 0 5888 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_70
timestamp 1729294469
transform 1 0 6992 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_82
timestamp 1729294469
transform 1 0 8096 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_94
timestamp 1729294469
transform 1 0 9200 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_102
timestamp 1729294469
transform 1 0 9936 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_112
timestamp 1729294469
transform 1 0 10856 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_124
timestamp 1729294469
transform 1 0 11960 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_132
timestamp 1729294469
transform 1 0 12696 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_157
timestamp 1729294469
transform 1 0 14996 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_167
timestamp 1729294469
transform 1 0 15916 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_171
timestamp 1729294469
transform 1 0 16284 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_186
timestamp 1729294469
transform 1 0 17664 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_192
timestamp 1729294469
transform 1 0 18216 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_207
timestamp 1729294469
transform 1 0 19596 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_215
timestamp 1729294469
transform 1 0 20332 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_242
timestamp 1729294469
transform 1 0 22816 0 1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1729294469
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1729294469
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_27
timestamp 1729294469
transform 1 0 3036 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_35
timestamp 1729294469
transform 1 0 3772 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_50
timestamp 1729294469
transform 1 0 5152 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_57
timestamp 1729294469
transform 1 0 5796 0 -1 10336
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_84
timestamp 1729294469
transform 1 0 8280 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_96
timestamp 1729294469
transform 1 0 9384 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_108
timestamp 1729294469
transform 1 0 10488 0 -1 10336
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1729294469
transform 1 0 10948 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_125
timestamp 1729294469
transform 1 0 12052 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_131
timestamp 1729294469
transform 1 0 12604 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_154
timestamp 1729294469
transform 1 0 14720 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_162
timestamp 1729294469
transform 1 0 15456 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_182
timestamp 1729294469
transform 1 0 17296 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_196
timestamp 1729294469
transform 1 0 18584 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_204
timestamp 1729294469
transform 1 0 19320 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_213
timestamp 1729294469
transform 1 0 20148 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_221
timestamp 1729294469
transform 1 0 20884 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_242
timestamp 1729294469
transform 1 0 22816 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1729294469
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1729294469
transform 1 0 1932 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1729294469
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1729294469
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_41
timestamp 1729294469
transform 1 0 4324 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_49
timestamp 1729294469
transform 1 0 5060 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_68
timestamp 1729294469
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_130
timestamp 1729294469
transform 1 0 12512 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_138
timestamp 1729294469
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_141
timestamp 1729294469
transform 1 0 13524 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_151
timestamp 1729294469
transform 1 0 14444 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_163
timestamp 1729294469
transform 1 0 15548 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_175
timestamp 1729294469
transform 1 0 16652 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_179
timestamp 1729294469
transform 1 0 17020 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_225
timestamp 1729294469
transform 1 0 21252 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_237
timestamp 1729294469
transform 1 0 22356 0 1 10336
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1729294469
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1729294469
transform 1 0 1932 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_27
timestamp 1729294469
transform 1 0 3036 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_45
timestamp 1729294469
transform 1 0 4692 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_53
timestamp 1729294469
transform 1 0 5428 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_66
timestamp 1729294469
transform 1 0 6624 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_78
timestamp 1729294469
transform 1 0 7728 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_84
timestamp 1729294469
transform 1 0 8280 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_96
timestamp 1729294469
transform 1 0 9384 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_104
timestamp 1729294469
transform 1 0 10120 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_113
timestamp 1729294469
transform 1 0 10948 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_123
timestamp 1729294469
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_135
timestamp 1729294469
transform 1 0 12972 0 -1 11424
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_146
timestamp 1729294469
transform 1 0 13984 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_158
timestamp 1729294469
transform 1 0 15088 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 1729294469
transform 1 0 16100 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_181
timestamp 1729294469
transform 1 0 17204 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_189
timestamp 1729294469
transform 1 0 17940 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_197
timestamp 1729294469
transform 1 0 18676 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_213
timestamp 1729294469
transform 1 0 20148 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1729294469
transform 1 0 21068 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_236
timestamp 1729294469
transform 1 0 22264 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_244
timestamp 1729294469
transform 1 0 23000 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1729294469
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1729294469
transform 1 0 1932 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1729294469
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_54
timestamp 1729294469
transform 1 0 5520 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_66
timestamp 1729294469
transform 1 0 6624 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_74
timestamp 1729294469
transform 1 0 7360 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1729294469
transform 1 0 8188 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_90
timestamp 1729294469
transform 1 0 8832 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_98
timestamp 1729294469
transform 1 0 9568 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_102
timestamp 1729294469
transform 1 0 9936 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_114
timestamp 1729294469
transform 1 0 11040 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_126
timestamp 1729294469
transform 1 0 12144 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_138
timestamp 1729294469
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_157
timestamp 1729294469
transform 1 0 14996 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_165
timestamp 1729294469
transform 1 0 15732 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_177
timestamp 1729294469
transform 1 0 16836 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_181
timestamp 1729294469
transform 1 0 17204 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_187
timestamp 1729294469
transform 1 0 17756 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1729294469
transform 1 0 18492 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_197
timestamp 1729294469
transform 1 0 18676 0 1 11424
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1729294469
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1729294469
transform 1 0 1932 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_36
timestamp 1729294469
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_53
timestamp 1729294469
transform 1 0 5428 0 -1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1729294469
transform 1 0 5796 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_69
timestamp 1729294469
transform 1 0 6900 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_76
timestamp 1729294469
transform 1 0 7544 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_80
timestamp 1729294469
transform 1 0 7912 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_89
timestamp 1729294469
transform 1 0 8740 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_95
timestamp 1729294469
transform 1 0 9292 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_109
timestamp 1729294469
transform 1 0 10580 0 -1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1729294469
transform 1 0 10948 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_125
timestamp 1729294469
transform 1 0 12052 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_131
timestamp 1729294469
transform 1 0 12604 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_135
timestamp 1729294469
transform 1 0 12972 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_143
timestamp 1729294469
transform 1 0 13708 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_151
timestamp 1729294469
transform 1 0 14444 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_169
timestamp 1729294469
transform 1 0 16100 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_184
timestamp 1729294469
transform 1 0 17480 0 -1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_202
timestamp 1729294469
transform 1 0 19136 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1729294469
transform 1 0 21068 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_225
timestamp 1729294469
transform 1 0 21252 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_238
timestamp 1729294469
transform 1 0 22448 0 -1 12512
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1729294469
transform 1 0 828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1729294469
transform 1 0 1932 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1729294469
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1729294469
transform 1 0 3220 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_41
timestamp 1729294469
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_52
timestamp 1729294469
transform 1 0 5336 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_64
timestamp 1729294469
transform 1 0 6440 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_78
timestamp 1729294469
transform 1 0 7728 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_85
timestamp 1729294469
transform 1 0 8372 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1729294469
transform 1 0 9476 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 1729294469
transform 1 0 10580 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1729294469
transform 1 0 13340 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_145
timestamp 1729294469
transform 1 0 13892 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_153
timestamp 1729294469
transform 1 0 14628 0 1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_165
timestamp 1729294469
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_177
timestamp 1729294469
transform 1 0 16836 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1729294469
transform 1 0 18492 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 1729294469
transform 1 0 18676 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_209
timestamp 1729294469
transform 1 0 19780 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_221
timestamp 1729294469
transform 1 0 20884 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_229
timestamp 1729294469
transform 1 0 21620 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_234
timestamp 1729294469
transform 1 0 22080 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_242
timestamp 1729294469
transform 1 0 22816 0 1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1729294469
transform 1 0 828 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_15
timestamp 1729294469
transform 1 0 1932 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_23
timestamp 1729294469
transform 1 0 2668 0 -1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_42
timestamp 1729294469
transform 1 0 4416 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_54
timestamp 1729294469
transform 1 0 5520 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_57
timestamp 1729294469
transform 1 0 5796 0 -1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_63
timestamp 1729294469
transform 1 0 6348 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_75
timestamp 1729294469
transform 1 0 7452 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_87
timestamp 1729294469
transform 1 0 8556 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_95
timestamp 1729294469
transform 1 0 9292 0 -1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1729294469
transform 1 0 10948 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_125
timestamp 1729294469
transform 1 0 12052 0 -1 13600
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_153
timestamp 1729294469
transform 1 0 14628 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_165
timestamp 1729294469
transform 1 0 15732 0 -1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1729294469
transform 1 0 16100 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_181
timestamp 1729294469
transform 1 0 17204 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_187
timestamp 1729294469
transform 1 0 17756 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_199
timestamp 1729294469
transform 1 0 18860 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_211
timestamp 1729294469
transform 1 0 19964 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1729294469
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_225
timestamp 1729294469
transform 1 0 21252 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_243
timestamp 1729294469
transform 1 0 22908 0 -1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1729294469
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_15
timestamp 1729294469
transform 1 0 1932 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_23
timestamp 1729294469
transform 1 0 2668 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_36
timestamp 1729294469
transform 1 0 3864 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_48
timestamp 1729294469
transform 1 0 4968 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_57
timestamp 1729294469
transform 1 0 5796 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_77
timestamp 1729294469
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_85
timestamp 1729294469
transform 1 0 8372 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_95
timestamp 1729294469
transform 1 0 9292 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_104
timestamp 1729294469
transform 1 0 10120 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_108
timestamp 1729294469
transform 1 0 10488 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_112
timestamp 1729294469
transform 1 0 10856 0 1 13600
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_127
timestamp 1729294469
transform 1 0 12236 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1729294469
transform 1 0 13340 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_148
timestamp 1729294469
transform 1 0 14168 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_192
timestamp 1729294469
transform 1 0 18216 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_211
timestamp 1729294469
transform 1 0 19964 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_224
timestamp 1729294469
transform 1 0 21160 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_243
timestamp 1729294469
transform 1 0 22908 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1729294469
transform 1 0 828 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_15
timestamp 1729294469
transform 1 0 1932 0 -1 14688
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_28
timestamp 1729294469
transform 1 0 3128 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_40
timestamp 1729294469
transform 1 0 4232 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_44
timestamp 1729294469
transform 1 0 4600 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1729294469
transform 1 0 5612 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_64
timestamp 1729294469
transform 1 0 6440 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_76
timestamp 1729294469
transform 1 0 7544 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_86
timestamp 1729294469
transform 1 0 8464 0 -1 14688
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_99
timestamp 1729294469
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1729294469
transform 1 0 10764 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1729294469
transform 1 0 10948 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1729294469
transform 1 0 12052 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 1729294469
transform 1 0 13156 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 1729294469
transform 1 0 14260 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_176
timestamp 1729294469
transform 1 0 16744 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_188
timestamp 1729294469
transform 1 0 17848 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_212
timestamp 1729294469
transform 1 0 20056 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_220
timestamp 1729294469
transform 1 0 20792 0 -1 14688
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1729294469
transform 1 0 21252 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_237
timestamp 1729294469
transform 1 0 22356 0 -1 14688
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1729294469
transform 1 0 828 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1729294469
transform 1 0 1932 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1729294469
transform 1 0 3036 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_29
timestamp 1729294469
transform 1 0 3220 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_51
timestamp 1729294469
transform 1 0 5244 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_60
timestamp 1729294469
transform 1 0 6072 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_72
timestamp 1729294469
transform 1 0 7176 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1729294469
transform 1 0 8372 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1729294469
transform 1 0 9476 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_109
timestamp 1729294469
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_118
timestamp 1729294469
transform 1 0 11408 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_126
timestamp 1729294469
transform 1 0 12144 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_146
timestamp 1729294469
transform 1 0 13984 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_158
timestamp 1729294469
transform 1 0 15088 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_166
timestamp 1729294469
transform 1 0 15824 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_178
timestamp 1729294469
transform 1 0 16928 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_190
timestamp 1729294469
transform 1 0 18032 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_200
timestamp 1729294469
transform 1 0 18952 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_208
timestamp 1729294469
transform 1 0 19688 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_215
timestamp 1729294469
transform 1 0 20332 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_221
timestamp 1729294469
transform 1 0 20884 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_229
timestamp 1729294469
transform 1 0 21620 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_236
timestamp 1729294469
transform 1 0 22264 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_244
timestamp 1729294469
transform 1 0 23000 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1729294469
transform 1 0 828 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_15
timestamp 1729294469
transform 1 0 1932 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_23
timestamp 1729294469
transform 1 0 2668 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_47
timestamp 1729294469
transform 1 0 4876 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1729294469
transform 1 0 5612 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1729294469
transform 1 0 5796 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_69
timestamp 1729294469
transform 1 0 6900 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_77
timestamp 1729294469
transform 1 0 7636 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_88
timestamp 1729294469
transform 1 0 8648 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_100
timestamp 1729294469
transform 1 0 9752 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_125
timestamp 1729294469
transform 1 0 12052 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_133
timestamp 1729294469
transform 1 0 12788 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_150
timestamp 1729294469
transform 1 0 14352 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1729294469
transform 1 0 15916 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1729294469
transform 1 0 16100 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_181
timestamp 1729294469
transform 1 0 17204 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_189
timestamp 1729294469
transform 1 0 17940 0 -1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_208
timestamp 1729294469
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_220
timestamp 1729294469
transform 1 0 20792 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_225
timestamp 1729294469
transform 1 0 21252 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_241
timestamp 1729294469
transform 1 0 22724 0 -1 15776
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1729294469
transform 1 0 828 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_15
timestamp 1729294469
transform 1 0 1932 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_41
timestamp 1729294469
transform 1 0 4324 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_49
timestamp 1729294469
transform 1 0 5060 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_65
timestamp 1729294469
transform 1 0 6532 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_69
timestamp 1729294469
transform 1 0 6900 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_103
timestamp 1729294469
transform 1 0 10028 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_119
timestamp 1729294469
transform 1 0 11500 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_131
timestamp 1729294469
transform 1 0 12604 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_146
timestamp 1729294469
transform 1 0 13984 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_154
timestamp 1729294469
transform 1 0 14720 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_160
timestamp 1729294469
transform 1 0 15272 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_184
timestamp 1729294469
transform 1 0 17480 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_188
timestamp 1729294469
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1729294469
transform 1 0 18492 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_208
timestamp 1729294469
transform 1 0 19688 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_220
timestamp 1729294469
transform 1 0 20792 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_226
timestamp 1729294469
transform 1 0 21344 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_235
timestamp 1729294469
transform 1 0 22172 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_243
timestamp 1729294469
transform 1 0 22908 0 1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1729294469
transform 1 0 828 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_15
timestamp 1729294469
transform 1 0 1932 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_23
timestamp 1729294469
transform 1 0 2668 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1729294469
transform 1 0 5612 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_57
timestamp 1729294469
transform 1 0 5796 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_78
timestamp 1729294469
transform 1 0 7728 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_82
timestamp 1729294469
transform 1 0 8096 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_88
timestamp 1729294469
transform 1 0 8648 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_100
timestamp 1729294469
transform 1 0 9752 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_104
timestamp 1729294469
transform 1 0 10120 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_134
timestamp 1729294469
transform 1 0 12880 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_142
timestamp 1729294469
transform 1 0 13616 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_147
timestamp 1729294469
transform 1 0 14076 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_155
timestamp 1729294469
transform 1 0 14812 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_177
timestamp 1729294469
transform 1 0 16836 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_213
timestamp 1729294469
transform 1 0 20148 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_221
timestamp 1729294469
transform 1 0 20884 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_225
timestamp 1729294469
transform 1 0 21252 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_243
timestamp 1729294469
transform 1 0 22908 0 -1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1729294469
transform 1 0 828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1729294469
transform 1 0 1932 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1729294469
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_29
timestamp 1729294469
transform 1 0 3220 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_33
timestamp 1729294469
transform 1 0 3588 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_39
timestamp 1729294469
transform 1 0 4140 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_51
timestamp 1729294469
transform 1 0 5244 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_57
timestamp 1729294469
transform 1 0 5796 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_61
timestamp 1729294469
transform 1 0 6164 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_73
timestamp 1729294469
transform 1 0 7268 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_81
timestamp 1729294469
transform 1 0 8004 0 1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_92
timestamp 1729294469
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_104
timestamp 1729294469
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_116
timestamp 1729294469
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_128
timestamp 1729294469
transform 1 0 12328 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_148
timestamp 1729294469
transform 1 0 14168 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_160
timestamp 1729294469
transform 1 0 15272 0 1 16864
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_169
timestamp 1729294469
transform 1 0 16100 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_181
timestamp 1729294469
transform 1 0 17204 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_187
timestamp 1729294469
transform 1 0 17756 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1729294469
transform 1 0 18492 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_204
timestamp 1729294469
transform 1 0 19320 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_232
timestamp 1729294469
transform 1 0 21896 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_244
timestamp 1729294469
transform 1 0 23000 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1729294469
transform 1 0 828 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1729294469
transform 1 0 1932 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_27
timestamp 1729294469
transform 1 0 3036 0 -1 17952
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_41
timestamp 1729294469
transform 1 0 4324 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_53
timestamp 1729294469
transform 1 0 5428 0 -1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1729294469
transform 1 0 5796 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1729294469
transform 1 0 6900 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 1729294469
transform 1 0 8004 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_93
timestamp 1729294469
transform 1 0 9108 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_108
timestamp 1729294469
transform 1 0 10488 0 -1 17952
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1729294469
transform 1 0 10948 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_125
timestamp 1729294469
transform 1 0 12052 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_133
timestamp 1729294469
transform 1 0 12788 0 -1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_154
timestamp 1729294469
transform 1 0 14720 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_166
timestamp 1729294469
transform 1 0 15824 0 -1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1729294469
transform 1 0 16100 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_181
timestamp 1729294469
transform 1 0 17204 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_185
timestamp 1729294469
transform 1 0 17572 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_189
timestamp 1729294469
transform 1 0 17940 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_201
timestamp 1729294469
transform 1 0 19044 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_213
timestamp 1729294469
transform 1 0 20148 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_221
timestamp 1729294469
transform 1 0 20884 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_225
timestamp 1729294469
transform 1 0 21252 0 -1 17952
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_233
timestamp 1729294469
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1729294469
transform 1 0 828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1729294469
transform 1 0 1932 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1729294469
transform 1 0 3036 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_29
timestamp 1729294469
transform 1 0 3220 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_37
timestamp 1729294469
transform 1 0 3956 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_54
timestamp 1729294469
transform 1 0 5520 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_66
timestamp 1729294469
transform 1 0 6624 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_72
timestamp 1729294469
transform 1 0 7176 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_79
timestamp 1729294469
transform 1 0 7820 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1729294469
transform 1 0 8188 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_85
timestamp 1729294469
transform 1 0 8372 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_90
timestamp 1729294469
transform 1 0 8832 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_124
timestamp 1729294469
transform 1 0 11960 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_138
timestamp 1729294469
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_148
timestamp 1729294469
transform 1 0 14168 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_156
timestamp 1729294469
transform 1 0 14904 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_174
timestamp 1729294469
transform 1 0 16560 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_180
timestamp 1729294469
transform 1 0 17112 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_186
timestamp 1729294469
transform 1 0 17664 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_194
timestamp 1729294469
transform 1 0 18400 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_197
timestamp 1729294469
transform 1 0 18676 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_205
timestamp 1729294469
transform 1 0 19412 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_213
timestamp 1729294469
transform 1 0 20148 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_224
timestamp 1729294469
transform 1 0 21160 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_228
timestamp 1729294469
transform 1 0 21528 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1729294469
transform 1 0 828 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_15
timestamp 1729294469
transform 1 0 1932 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_23
timestamp 1729294469
transform 1 0 2668 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_30
timestamp 1729294469
transform 1 0 3312 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_78
timestamp 1729294469
transform 1 0 7728 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1729294469
transform 1 0 10764 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_113
timestamp 1729294469
transform 1 0 10948 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_121
timestamp 1729294469
transform 1 0 11684 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_140
timestamp 1729294469
transform 1 0 13432 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_148
timestamp 1729294469
transform 1 0 14168 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_158
timestamp 1729294469
transform 1 0 15088 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_166
timestamp 1729294469
transform 1 0 15824 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_169
timestamp 1729294469
transform 1 0 16100 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_178
timestamp 1729294469
transform 1 0 16928 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_184
timestamp 1729294469
transform 1 0 17480 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_189
timestamp 1729294469
transform 1 0 17940 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_196
timestamp 1729294469
transform 1 0 18584 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_215
timestamp 1729294469
transform 1 0 20332 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1729294469
transform 1 0 828 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_15
timestamp 1729294469
transform 1 0 1932 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_21
timestamp 1729294469
transform 1 0 2484 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_41
timestamp 1729294469
transform 1 0 4324 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_45
timestamp 1729294469
transform 1 0 4692 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_53
timestamp 1729294469
transform 1 0 5428 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_77
timestamp 1729294469
transform 1 0 7636 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1729294469
transform 1 0 8188 0 1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_85
timestamp 1729294469
transform 1 0 8372 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_119
timestamp 1729294469
transform 1 0 11500 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_129
timestamp 1729294469
transform 1 0 12420 0 1 19040
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_141
timestamp 1729294469
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_153
timestamp 1729294469
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_165
timestamp 1729294469
transform 1 0 15732 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_181
timestamp 1729294469
transform 1 0 17204 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_194
timestamp 1729294469
transform 1 0 18400 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_210
timestamp 1729294469
transform 1 0 19872 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_214
timestamp 1729294469
transform 1 0 20240 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_230
timestamp 1729294469
transform 1 0 21712 0 1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1729294469
transform 1 0 828 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_15
timestamp 1729294469
transform 1 0 1932 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_33
timestamp 1729294469
transform 1 0 3588 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_44
timestamp 1729294469
transform 1 0 4600 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_48
timestamp 1729294469
transform 1 0 4968 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1729294469
transform 1 0 5612 0 -1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1729294469
transform 1 0 5796 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_69
timestamp 1729294469
transform 1 0 6900 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_106
timestamp 1729294469
transform 1 0 10304 0 -1 20128
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_120
timestamp 1729294469
transform 1 0 11592 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_132
timestamp 1729294469
transform 1 0 12696 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_144
timestamp 1729294469
transform 1 0 13800 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_156
timestamp 1729294469
transform 1 0 14904 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 1729294469
transform 1 0 16100 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_181
timestamp 1729294469
transform 1 0 17204 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_193
timestamp 1729294469
transform 1 0 18308 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_203
timestamp 1729294469
transform 1 0 19228 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_211
timestamp 1729294469
transform 1 0 19964 0 -1 20128
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_233
timestamp 1729294469
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1729294469
transform 1 0 828 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1729294469
transform 1 0 1932 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1729294469
transform 1 0 3036 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_29
timestamp 1729294469
transform 1 0 3220 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_37
timestamp 1729294469
transform 1 0 3956 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_49
timestamp 1729294469
transform 1 0 5060 0 1 20128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_57
timestamp 1729294469
transform 1 0 5796 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_69
timestamp 1729294469
transform 1 0 6900 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_81
timestamp 1729294469
transform 1 0 8004 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_85
timestamp 1729294469
transform 1 0 8372 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_93
timestamp 1729294469
transform 1 0 9108 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_97
timestamp 1729294469
transform 1 0 9476 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_109
timestamp 1729294469
transform 1 0 10580 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_121
timestamp 1729294469
transform 1 0 11684 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_133
timestamp 1729294469
transform 1 0 12788 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1729294469
transform 1 0 13340 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_141
timestamp 1729294469
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_153
timestamp 1729294469
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_165
timestamp 1729294469
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_177
timestamp 1729294469
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_189
timestamp 1729294469
transform 1 0 17940 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 1729294469
transform 1 0 18492 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_197
timestamp 1729294469
transform 1 0 18676 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_208
timestamp 1729294469
transform 1 0 19688 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_216
timestamp 1729294469
transform 1 0 20424 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_231
timestamp 1729294469
transform 1 0 21804 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_243
timestamp 1729294469
transform 1 0 22908 0 1 20128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1729294469
transform 1 0 828 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1729294469
transform 1 0 1932 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_27
timestamp 1729294469
transform 1 0 3036 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_33
timestamp 1729294469
transform 1 0 3588 0 -1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1729294469
transform 1 0 5796 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_69
timestamp 1729294469
transform 1 0 6900 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_79
timestamp 1729294469
transform 1 0 7820 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_90
timestamp 1729294469
transform 1 0 8832 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_97
timestamp 1729294469
transform 1 0 9476 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_104
timestamp 1729294469
transform 1 0 10120 0 -1 21216
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 1729294469
transform 1 0 10948 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_125
timestamp 1729294469
transform 1 0 12052 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_148
timestamp 1729294469
transform 1 0 14168 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_157
timestamp 1729294469
transform 1 0 14996 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_164
timestamp 1729294469
transform 1 0 15640 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_169
timestamp 1729294469
transform 1 0 16100 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_175
timestamp 1729294469
transform 1 0 16652 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_180
timestamp 1729294469
transform 1 0 17112 0 -1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_188
timestamp 1729294469
transform 1 0 17848 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_200
timestamp 1729294469
transform 1 0 18952 0 -1 21216
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_209
timestamp 1729294469
transform 1 0 19780 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_221
timestamp 1729294469
transform 1 0 20884 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_238
timestamp 1729294469
transform 1 0 22448 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_244
timestamp 1729294469
transform 1 0 23000 0 -1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1729294469
transform 1 0 828 0 1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1729294469
transform 1 0 1932 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1729294469
transform 1 0 3036 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_29
timestamp 1729294469
transform 1 0 3220 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_71
timestamp 1729294469
transform 1 0 7084 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_115
timestamp 1729294469
transform 1 0 11132 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_166
timestamp 1729294469
transform 1 0 15824 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_173
timestamp 1729294469
transform 1 0 16468 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 1729294469
transform 1 0 18492 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_197
timestamp 1729294469
transform 1 0 18676 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_205
timestamp 1729294469
transform 1 0 19412 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_211
timestamp 1729294469
transform 1 0 19964 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_215
timestamp 1729294469
transform 1 0 20332 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_234
timestamp 1729294469
transform 1 0 22080 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_242
timestamp 1729294469
transform 1 0 22816 0 1 21216
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1729294469
transform 1 0 828 0 -1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1729294469
transform 1 0 1932 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_27
timestamp 1729294469
transform 1 0 3036 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_33
timestamp 1729294469
transform 1 0 3588 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_60
timestamp 1729294469
transform 1 0 6072 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_92
timestamp 1729294469
transform 1 0 9016 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_148
timestamp 1729294469
transform 1 0 14168 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_152
timestamp 1729294469
transform 1 0 14536 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_165
timestamp 1729294469
transform 1 0 15732 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_184
timestamp 1729294469
transform 1 0 17480 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_189
timestamp 1729294469
transform 1 0 17940 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_206
timestamp 1729294469
transform 1 0 19504 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_242
timestamp 1729294469
transform 1 0 22816 0 -1 22304
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1729294469
transform 1 0 828 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_15
timestamp 1729294469
transform 1 0 1932 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_23
timestamp 1729294469
transform 1 0 2668 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_29
timestamp 1729294469
transform 1 0 3220 0 1 22304
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_61
timestamp 1729294469
transform 1 0 6164 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_80
timestamp 1729294469
transform 1 0 7912 0 1 22304
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_90
timestamp 1729294469
transform 1 0 8832 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_102
timestamp 1729294469
transform 1 0 9936 0 1 22304
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_109
timestamp 1729294469
transform 1 0 10580 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_121
timestamp 1729294469
transform 1 0 11684 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_126
timestamp 1729294469
transform 1 0 12144 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_137
timestamp 1729294469
transform 1 0 13156 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_141
timestamp 1729294469
transform 1 0 13524 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_150
timestamp 1729294469
transform 1 0 14352 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_176
timestamp 1729294469
transform 1 0 16744 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_182
timestamp 1729294469
transform 1 0 17296 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1729294469
transform 1 0 18492 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_210
timestamp 1729294469
transform 1 0 19872 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_214
timestamp 1729294469
transform 1 0 20240 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_219
timestamp 1729294469
transform 1 0 20700 0 1 22304
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_233
timestamp 1729294469
transform 1 0 21988 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_3
timestamp 1729294469
transform 1 0 828 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_11
timestamp 1729294469
transform 1 0 1564 0 -1 23392
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_16
timestamp 1729294469
transform 1 0 2024 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_29
timestamp 1729294469
transform 1 0 3220 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_36
timestamp 1729294469
transform 1 0 3864 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_53
timestamp 1729294469
transform 1 0 5428 0 -1 23392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1729294469
transform 1 0 5796 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_69
timestamp 1729294469
transform 1 0 6900 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_80
timestamp 1729294469
transform 1 0 7912 0 -1 23392
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_85
timestamp 1729294469
transform 1 0 8372 0 -1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_97
timestamp 1729294469
transform 1 0 9476 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_109
timestamp 1729294469
transform 1 0 10580 0 -1 23392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_119
timestamp 1729294469
transform 1 0 11500 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_131
timestamp 1729294469
transform 1 0 12604 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_139
timestamp 1729294469
transform 1 0 13340 0 -1 23392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_147
timestamp 1729294469
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_159
timestamp 1729294469
transform 1 0 15180 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 1729294469
transform 1 0 15916 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_169
timestamp 1729294469
transform 1 0 16100 0 -1 23392
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_176
timestamp 1729294469
transform 1 0 16744 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_188
timestamp 1729294469
transform 1 0 17848 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_192
timestamp 1729294469
transform 1 0 18216 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_197
timestamp 1729294469
transform 1 0 18676 0 -1 23392
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_211
timestamp 1729294469
transform 1 0 19964 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 1729294469
transform 1 0 21068 0 -1 23392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 1729294469
transform 1 0 21252 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_243
timestamp 1729294469
transform 1 0 22908 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1729294469
transform -1 0 23092 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1729294469
transform 1 0 22816 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1729294469
transform 1 0 1748 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1729294469
transform -1 0 5428 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1729294469
transform -1 0 7912 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input6
timestamp 1729294469
transform 1 0 10948 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input7
timestamp 1729294469
transform 1 0 13524 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1729294469
transform 1 0 16468 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input9
timestamp 1729294469
transform 1 0 19412 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input10
timestamp 1729294469
transform 1 0 22356 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_42
timestamp 1729294469
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1729294469
transform -1 0 23368 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_43
timestamp 1729294469
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1729294469
transform -1 0 23368 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_44
timestamp 1729294469
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1729294469
transform -1 0 23368 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_45
timestamp 1729294469
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1729294469
transform -1 0 23368 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_46
timestamp 1729294469
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1729294469
transform -1 0 23368 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_47
timestamp 1729294469
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1729294469
transform -1 0 23368 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_48
timestamp 1729294469
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1729294469
transform -1 0 23368 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_49
timestamp 1729294469
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1729294469
transform -1 0 23368 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_50
timestamp 1729294469
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1729294469
transform -1 0 23368 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_51
timestamp 1729294469
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1729294469
transform -1 0 23368 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_52
timestamp 1729294469
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1729294469
transform -1 0 23368 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_53
timestamp 1729294469
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1729294469
transform -1 0 23368 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_54
timestamp 1729294469
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1729294469
transform -1 0 23368 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_55
timestamp 1729294469
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1729294469
transform -1 0 23368 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_56
timestamp 1729294469
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1729294469
transform -1 0 23368 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_57
timestamp 1729294469
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1729294469
transform -1 0 23368 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_58
timestamp 1729294469
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1729294469
transform -1 0 23368 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_59
timestamp 1729294469
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1729294469
transform -1 0 23368 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_60
timestamp 1729294469
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1729294469
transform -1 0 23368 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_61
timestamp 1729294469
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1729294469
transform -1 0 23368 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_62
timestamp 1729294469
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1729294469
transform -1 0 23368 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_63
timestamp 1729294469
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1729294469
transform -1 0 23368 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_64
timestamp 1729294469
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1729294469
transform -1 0 23368 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_65
timestamp 1729294469
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1729294469
transform -1 0 23368 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_66
timestamp 1729294469
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1729294469
transform -1 0 23368 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_67
timestamp 1729294469
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1729294469
transform -1 0 23368 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_68
timestamp 1729294469
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1729294469
transform -1 0 23368 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_69
timestamp 1729294469
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1729294469
transform -1 0 23368 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_70
timestamp 1729294469
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1729294469
transform -1 0 23368 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_71
timestamp 1729294469
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1729294469
transform -1 0 23368 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_72
timestamp 1729294469
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1729294469
transform -1 0 23368 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_73
timestamp 1729294469
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1729294469
transform -1 0 23368 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_74
timestamp 1729294469
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1729294469
transform -1 0 23368 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_75
timestamp 1729294469
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1729294469
transform -1 0 23368 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_76
timestamp 1729294469
transform 1 0 552 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1729294469
transform -1 0 23368 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_77
timestamp 1729294469
transform 1 0 552 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1729294469
transform -1 0 23368 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_78
timestamp 1729294469
transform 1 0 552 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1729294469
transform -1 0 23368 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_79
timestamp 1729294469
transform 1 0 552 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1729294469
transform -1 0 23368 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_80
timestamp 1729294469
transform 1 0 552 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1729294469
transform -1 0 23368 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_81
timestamp 1729294469
transform 1 0 552 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1729294469
transform -1 0 23368 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_82
timestamp 1729294469
transform 1 0 552 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1729294469
transform -1 0 23368 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_83
timestamp 1729294469
transform 1 0 552 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1729294469
transform -1 0 23368 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_84
timestamp 1729294469
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_85
timestamp 1729294469
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_86
timestamp 1729294469
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_87
timestamp 1729294469
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_88
timestamp 1729294469
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_89
timestamp 1729294469
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_90
timestamp 1729294469
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_91
timestamp 1729294469
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_92
timestamp 1729294469
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_93
timestamp 1729294469
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_94
timestamp 1729294469
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_95
timestamp 1729294469
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_96
timestamp 1729294469
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_97
timestamp 1729294469
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_98
timestamp 1729294469
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_99
timestamp 1729294469
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_100
timestamp 1729294469
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_101
timestamp 1729294469
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_102
timestamp 1729294469
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_103
timestamp 1729294469
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_104
timestamp 1729294469
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_105
timestamp 1729294469
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_106
timestamp 1729294469
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_107
timestamp 1729294469
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_108
timestamp 1729294469
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_109
timestamp 1729294469
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_110
timestamp 1729294469
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_111
timestamp 1729294469
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_112
timestamp 1729294469
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_113
timestamp 1729294469
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_114
timestamp 1729294469
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_115
timestamp 1729294469
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_116
timestamp 1729294469
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_117
timestamp 1729294469
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_118
timestamp 1729294469
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_119
timestamp 1729294469
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_120
timestamp 1729294469
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_121
timestamp 1729294469
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_122
timestamp 1729294469
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_123
timestamp 1729294469
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_124
timestamp 1729294469
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_125
timestamp 1729294469
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_126
timestamp 1729294469
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_127
timestamp 1729294469
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_128
timestamp 1729294469
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_129
timestamp 1729294469
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_130
timestamp 1729294469
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_131
timestamp 1729294469
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_132
timestamp 1729294469
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_133
timestamp 1729294469
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_134
timestamp 1729294469
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_135
timestamp 1729294469
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_136
timestamp 1729294469
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_137
timestamp 1729294469
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_138
timestamp 1729294469
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_139
timestamp 1729294469
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_140
timestamp 1729294469
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_141
timestamp 1729294469
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_142
timestamp 1729294469
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_143
timestamp 1729294469
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_144
timestamp 1729294469
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_145
timestamp 1729294469
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_146
timestamp 1729294469
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_147
timestamp 1729294469
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_148
timestamp 1729294469
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_149
timestamp 1729294469
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_150
timestamp 1729294469
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_151
timestamp 1729294469
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_152
timestamp 1729294469
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_153
timestamp 1729294469
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_154
timestamp 1729294469
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_155
timestamp 1729294469
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_156
timestamp 1729294469
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_157
timestamp 1729294469
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_158
timestamp 1729294469
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_159
timestamp 1729294469
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_160
timestamp 1729294469
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_161
timestamp 1729294469
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_162
timestamp 1729294469
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_163
timestamp 1729294469
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_164
timestamp 1729294469
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_165
timestamp 1729294469
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_166
timestamp 1729294469
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_167
timestamp 1729294469
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_168
timestamp 1729294469
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_169
timestamp 1729294469
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_170
timestamp 1729294469
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_171
timestamp 1729294469
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_172
timestamp 1729294469
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_173
timestamp 1729294469
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_174
timestamp 1729294469
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_175
timestamp 1729294469
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_176
timestamp 1729294469
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_177
timestamp 1729294469
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_178
timestamp 1729294469
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_179
timestamp 1729294469
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_180
timestamp 1729294469
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_181
timestamp 1729294469
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_182
timestamp 1729294469
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_183
timestamp 1729294469
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_184
timestamp 1729294469
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_185
timestamp 1729294469
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_186
timestamp 1729294469
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_187
timestamp 1729294469
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_188
timestamp 1729294469
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_189
timestamp 1729294469
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_190
timestamp 1729294469
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_191
timestamp 1729294469
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_192
timestamp 1729294469
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_193
timestamp 1729294469
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_194
timestamp 1729294469
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_195
timestamp 1729294469
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_196
timestamp 1729294469
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_197
timestamp 1729294469
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_198
timestamp 1729294469
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_199
timestamp 1729294469
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_200
timestamp 1729294469
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_201
timestamp 1729294469
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_202
timestamp 1729294469
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_203
timestamp 1729294469
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_204
timestamp 1729294469
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_205
timestamp 1729294469
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_206
timestamp 1729294469
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_207
timestamp 1729294469
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_208
timestamp 1729294469
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_209
timestamp 1729294469
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_210
timestamp 1729294469
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_211
timestamp 1729294469
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_212
timestamp 1729294469
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_213
timestamp 1729294469
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_214
timestamp 1729294469
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_215
timestamp 1729294469
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_216
timestamp 1729294469
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_217
timestamp 1729294469
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_218
timestamp 1729294469
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_219
timestamp 1729294469
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_220
timestamp 1729294469
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_221
timestamp 1729294469
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_222
timestamp 1729294469
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_223
timestamp 1729294469
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_224
timestamp 1729294469
transform 1 0 3128 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_225
timestamp 1729294469
transform 1 0 8280 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_226
timestamp 1729294469
transform 1 0 13432 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_227
timestamp 1729294469
transform 1 0 18584 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_228
timestamp 1729294469
transform 1 0 5704 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_229
timestamp 1729294469
transform 1 0 10856 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_230
timestamp 1729294469
transform 1 0 16008 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_231
timestamp 1729294469
transform 1 0 21160 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_232
timestamp 1729294469
transform 1 0 3128 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_233
timestamp 1729294469
transform 1 0 8280 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_234
timestamp 1729294469
transform 1 0 13432 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_235
timestamp 1729294469
transform 1 0 18584 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_236
timestamp 1729294469
transform 1 0 5704 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_237
timestamp 1729294469
transform 1 0 10856 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_238
timestamp 1729294469
transform 1 0 16008 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_239
timestamp 1729294469
transform 1 0 21160 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_240
timestamp 1729294469
transform 1 0 3128 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_241
timestamp 1729294469
transform 1 0 8280 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_242
timestamp 1729294469
transform 1 0 13432 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_243
timestamp 1729294469
transform 1 0 18584 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_244
timestamp 1729294469
transform 1 0 5704 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_245
timestamp 1729294469
transform 1 0 10856 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_246
timestamp 1729294469
transform 1 0 16008 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_247
timestamp 1729294469
transform 1 0 21160 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_248
timestamp 1729294469
transform 1 0 3128 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_249
timestamp 1729294469
transform 1 0 8280 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_250
timestamp 1729294469
transform 1 0 13432 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_251
timestamp 1729294469
transform 1 0 18584 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_252
timestamp 1729294469
transform 1 0 3128 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_253
timestamp 1729294469
transform 1 0 5704 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_254
timestamp 1729294469
transform 1 0 8280 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_255
timestamp 1729294469
transform 1 0 10856 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_256
timestamp 1729294469
transform 1 0 13432 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_257
timestamp 1729294469
transform 1 0 16008 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_258
timestamp 1729294469
transform 1 0 18584 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_259
timestamp 1729294469
transform 1 0 21160 0 -1 23392
box -38 -48 130 592
<< labels >>
rlabel metal1 s 11960 23392 11960 23392 4 VGND
rlabel metal1 s 11960 22848 11960 22848 4 VPWR
rlabel metal2 s 4374 11662 4374 11662 4 _0000_
rlabel metal1 s 3960 13430 3960 13430 4 _0001_
rlabel metal1 s 4135 11254 4135 11254 4 _0002_
rlabel metal2 s 4273 12342 4273 12342 4 _0003_
rlabel metal2 s 5653 10574 5653 10574 4 _0004_
rlabel metal2 s 7038 10302 7038 10302 4 _0005_
rlabel metal1 s 8229 9078 8229 9078 4 _0006_
rlabel metal1 s 9885 9078 9885 9078 4 _0007_
rlabel metal1 s 10161 10574 10161 10574 4 _0008_
rlabel metal1 s 11495 10574 11495 10574 4 _0009_
rlabel metal1 s 13896 11662 13896 11662 4 _0010_
rlabel metal1 s 14045 10166 14045 10166 4 _0011_
rlabel metal2 s 13841 9486 13841 9486 4 _0012_
rlabel metal1 s 14899 12342 14899 12342 4 _0013_
rlabel metal1 s 15492 13838 15492 13838 4 _0014_
rlabel metal1 s 16964 13838 16964 13838 4 _0015_
rlabel metal2 s 18533 15538 18533 15538 4 _0016_
rlabel metal2 s 19274 16422 19274 16422 4 _0017_
rlabel metal1 s 19223 18870 19223 18870 4 _0018_
rlabel metal1 s 20546 17034 20546 17034 4 _0019_
rlabel metal1 s 21840 18190 21840 18190 4 _0020_
rlabel metal2 s 21666 19006 21666 19006 4 _0021_
rlabel metal1 s 1876 4046 1876 4046 4 _0022_
rlabel metal2 s 4365 4046 4365 4046 4 _0023_
rlabel metal2 s 3537 3638 3537 3638 4 _0024_
rlabel metal1 s 2606 4726 2606 4726 4 _0025_
rlabel metal2 s 2162 7106 2162 7106 4 _0026_
rlabel metal1 s 3128 6970 3128 6970 4 _0027_
rlabel metal2 s 4830 6630 4830 6630 4 _0028_
rlabel metal1 s 5648 5134 5648 5134 4 _0029_
rlabel metal2 s 6389 5746 6389 5746 4 _0030_
rlabel metal1 s 8280 5338 8280 5338 4 _0031_
rlabel metal2 s 8965 4726 8965 4726 4 _0032_
rlabel metal2 s 10166 4930 10166 4930 4 _0033_
rlabel metal2 s 12102 5134 12102 5134 4 _0034_
rlabel metal1 s 13002 4726 13002 4726 4 _0035_
rlabel metal2 s 13841 5134 13841 5134 4 _0036_
rlabel metal1 s 15828 5134 15828 5134 4 _0037_
rlabel metal2 s 16422 6630 16422 6630 4 _0038_
rlabel metal1 s 15952 8398 15952 8398 4 _0039_
rlabel metal2 s 17530 9010 17530 9010 4 _0040_
rlabel metal1 s 19232 9078 19232 9078 4 _0041_
rlabel metal1 s 18507 10506 18507 10506 4 _0042_
rlabel metal2 s 20102 10370 20102 10370 4 _0043_
rlabel metal1 s 21026 11662 21026 11662 4 _0044_
rlabel metal2 s 21850 11458 21850 11458 4 _0045_
rlabel metal1 s 21466 9418 21466 9418 4 _0046_
rlabel metal1 s 21344 8602 21344 8602 4 _0047_
rlabel metal1 s 21650 6902 21650 6902 4 _0048_
rlabel metal1 s 21558 6154 21558 6154 4 _0049_
rlabel metal2 s 20005 4726 20005 4726 4 _0050_
rlabel metal1 s 18860 5338 18860 5338 4 _0051_
rlabel metal1 s 18676 6426 18676 6426 4 _0052_
rlabel metal2 s 18814 7718 18814 7718 4 _0053_
rlabel metal2 s 21753 16626 21753 16626 4 _0054_
rlabel metal2 s 22862 17544 22862 17544 4 _0055_
rlabel metal2 s 21022 19142 21022 19142 4 _0056_
rlabel metal2 s 3818 15742 3818 15742 4 _0057_
rlabel metal2 s 3542 16966 3542 16966 4 _0058_
rlabel metal1 s 6716 21318 6716 21318 4 _0059_
rlabel metal1 s 21298 21862 21298 21862 4 _0060_
rlabel metal2 s 5474 9860 5474 9860 4 _0061_
rlabel metal1 s 5888 8602 5888 8602 4 _0062_
rlabel metal1 s 8372 7854 8372 7854 4 _0063_
rlabel metal1 s 10626 8364 10626 8364 4 _0064_
rlabel metal1 s 11224 7854 11224 7854 4 _0065_
rlabel metal2 s 14122 8704 14122 8704 4 _0066_
rlabel metal1 s 13478 8466 13478 8466 4 _0067_
rlabel metal2 s 15686 9248 15686 9248 4 _0068_
rlabel metal1 s 17296 13362 17296 13362 4 _0069_
rlabel metal1 s 17756 12954 17756 12954 4 _0070_
rlabel metal1 s 20010 14382 20010 14382 4 _0071_
rlabel metal1 s 22218 15572 22218 15572 4 _0072_
rlabel metal2 s 22494 13022 22494 13022 4 _0073_
rlabel metal2 s 22862 10574 22862 10574 4 _0074_
rlabel metal1 s 3036 14586 3036 14586 4 _0075_
rlabel metal1 s 3174 13838 3174 13838 4 _0076_
rlabel metal2 s 3634 19108 3634 19108 4 _0077_
rlabel metal1 s 3358 19414 3358 19414 4 _0078_
rlabel metal1 s 3266 19346 3266 19346 4 _0079_
rlabel metal1 s 5060 11730 5060 11730 4 _0080_
rlabel metal1 s 3818 15674 3818 15674 4 _0081_
rlabel metal2 s 5842 22576 5842 22576 4 _0082_
rlabel metal1 s 4922 12614 4922 12614 4 _0083_
rlabel metal1 s 7406 18802 7406 18802 4 _0084_
rlabel metal1 s 9154 20366 9154 20366 4 _0085_
rlabel metal2 s 8235 21386 8235 21386 4 _0086_
rlabel metal1 s 6256 11322 6256 11322 4 _0087_
rlabel metal1 s 4830 22984 4830 22984 4 _0088_
rlabel metal1 s 4922 22678 4922 22678 4 _0089_
rlabel metal1 s 5612 21454 5612 21454 4 _0090_
rlabel metal1 s 7084 22134 7084 22134 4 _0091_
rlabel metal1 s 7314 12716 7314 12716 4 _0092_
rlabel metal1 s 8096 22474 8096 22474 4 _0093_
rlabel metal1 s 8648 22542 8648 22542 4 _0094_
rlabel metal2 s 5290 20468 5290 20468 4 _0095_
rlabel metal2 s 5014 16864 5014 16864 4 _0096_
rlabel metal2 s 3174 17136 3174 17136 4 _0097_
rlabel metal2 s 5106 17986 5106 17986 4 _0098_
rlabel metal2 s 6302 18768 6302 18768 4 _0099_
rlabel metal1 s 7360 19346 7360 19346 4 _0100_
rlabel metal1 s 8004 16694 8004 16694 4 _0101_
rlabel metal2 s 7590 18938 7590 18938 4 _0102_
rlabel metal1 s 8326 16422 8326 16422 4 _0103_
rlabel metal2 s 6946 15742 6946 15742 4 _0104_
rlabel metal1 s 8280 11594 8280 11594 4 _0105_
rlabel metal1 s 7268 12274 7268 12274 4 _0106_
rlabel metal1 s 7452 12274 7452 12274 4 _0107_
rlabel metal1 s 8050 12240 8050 12240 4 _0108_
rlabel metal1 s 8418 10540 8418 10540 4 _0109_
rlabel metal2 s 7590 11186 7590 11186 4 _0110_
rlabel metal2 s 10718 20060 10718 20060 4 _0111_
rlabel metal1 s 9154 14450 9154 14450 4 _0112_
rlabel metal1 s 8418 18802 8418 18802 4 _0113_
rlabel metal1 s 9154 18122 9154 18122 4 _0114_
rlabel metal1 s 3864 16626 3864 16626 4 _0115_
rlabel metal1 s 5934 16626 5934 16626 4 _0116_
rlabel metal2 s 6486 15810 6486 15810 4 _0117_
rlabel metal1 s 7314 15402 7314 15402 4 _0118_
rlabel metal2 s 8878 16558 8878 16558 4 _0119_
rlabel metal1 s 8280 16150 8280 16150 4 _0120_
rlabel metal1 s 8648 12274 8648 12274 4 _0121_
rlabel metal1 s 8648 12342 8648 12342 4 _0122_
rlabel metal2 s 8418 11866 8418 11866 4 _0123_
rlabel metal1 s 8510 11186 8510 11186 4 _0124_
rlabel metal2 s 8050 11356 8050 11356 4 _0125_
rlabel metal1 s 8326 10778 8326 10778 4 _0126_
rlabel metal2 s 8878 9996 8878 9996 4 _0127_
rlabel metal1 s 7176 13362 7176 13362 4 _0128_
rlabel metal1 s 5750 19380 5750 19380 4 _0129_
rlabel metal1 s 3542 15436 3542 15436 4 _0130_
rlabel metal2 s 5198 14620 5198 14620 4 _0131_
rlabel metal1 s 4232 16626 4232 16626 4 _0132_
rlabel metal1 s 5704 17102 5704 17102 4 _0133_
rlabel metal1 s 6026 13430 6026 13430 4 _0134_
rlabel metal2 s 6026 14110 6026 14110 4 _0135_
rlabel metal1 s 7789 13838 7789 13838 4 _0136_
rlabel metal1 s 8280 14382 8280 14382 4 _0137_
rlabel metal2 s 9522 13736 9522 13736 4 _0138_
rlabel metal2 s 8970 14076 8970 14076 4 _0139_
rlabel metal2 s 9706 13736 9706 13736 4 _0140_
rlabel metal1 s 8602 12750 8602 12750 4 _0141_
rlabel metal1 s 9798 12376 9798 12376 4 _0142_
rlabel metal2 s 9338 11866 9338 11866 4 _0143_
rlabel metal2 s 9154 11050 9154 11050 4 _0144_
rlabel metal1 s 8970 10642 8970 10642 4 _0145_
rlabel metal2 s 10534 9996 10534 9996 4 _0146_
rlabel metal2 s 15318 18564 15318 18564 4 _0147_
rlabel metal2 s 3358 18768 3358 18768 4 _0148_
rlabel metal2 s 7222 20859 7222 20859 4 _0149_
rlabel metal2 s 4186 15385 4186 15385 4 _0150_
rlabel metal2 s 4278 15164 4278 15164 4 _0151_
rlabel metal1 s 4968 14586 4968 14586 4 _0152_
rlabel metal1 s 5842 15028 5842 15028 4 _0153_
rlabel metal2 s 6762 14042 6762 14042 4 _0154_
rlabel metal2 s 6670 13566 6670 13566 4 _0155_
rlabel metal1 s 11362 13906 11362 13906 4 _0156_
rlabel metal1 s 10212 13838 10212 13838 4 _0157_
rlabel metal1 s 11362 14042 11362 14042 4 _0158_
rlabel metal2 s 10258 13532 10258 13532 4 _0159_
rlabel metal1 s 10028 11662 10028 11662 4 _0160_
rlabel metal1 s 10304 12274 10304 12274 4 _0161_
rlabel metal2 s 12466 12852 12466 12852 4 _0162_
rlabel metal1 s 10028 12070 10028 12070 4 _0163_
rlabel metal1 s 9614 12240 9614 12240 4 _0164_
rlabel metal1 s 10442 11730 10442 11730 4 _0165_
rlabel metal2 s 10718 11934 10718 11934 4 _0166_
rlabel metal1 s 10626 11628 10626 11628 4 _0167_
rlabel metal1 s 10856 11322 10856 11322 4 _0168_
rlabel metal1 s 16192 22542 16192 22542 4 _0169_
rlabel metal1 s 15916 22066 15916 22066 4 _0170_
rlabel metal1 s 15226 21998 15226 21998 4 _0171_
rlabel metal3 s 10350 22389 10350 22389 4 _0172_
rlabel metal1 s 16238 21352 16238 21352 4 _0173_
rlabel metal1 s 7774 22542 7774 22542 4 _0174_
rlabel metal1 s 7314 22406 7314 22406 4 _0175_
rlabel metal1 s 7774 21590 7774 21590 4 _0176_
rlabel metal1 s 10488 22474 10488 22474 4 _0177_
rlabel metal1 s 10442 22542 10442 22542 4 _0178_
rlabel metal2 s 10258 21692 10258 21692 4 _0179_
rlabel metal2 s 11362 18462 11362 18462 4 _0180_
rlabel metal2 s 11270 15300 11270 15300 4 _0181_
rlabel metal2 s 11638 15810 11638 15810 4 _0182_
rlabel metal2 s 10994 15742 10994 15742 4 _0183_
rlabel metal2 s 11546 14314 11546 14314 4 _0184_
rlabel metal1 s 13386 13294 13386 13294 4 _0185_
rlabel metal2 s 12742 13532 12742 13532 4 _0186_
rlabel metal2 s 13294 13634 13294 13634 4 _0187_
rlabel metal1 s 12604 12614 12604 12614 4 _0188_
rlabel metal2 s 11730 11900 11730 11900 4 _0189_
rlabel metal2 s 13570 11764 13570 11764 4 _0190_
rlabel metal1 s 13294 20944 13294 20944 4 _0191_
rlabel metal1 s 18584 22406 18584 22406 4 _0192_
rlabel metal1 s 18078 22066 18078 22066 4 _0193_
rlabel metal2 s 18354 22780 18354 22780 4 _0194_
rlabel metal2 s 19458 21692 19458 21692 4 _0195_
rlabel metal3 s 7314 21845 7314 21845 4 _0196_
rlabel metal2 s 11822 22338 11822 22338 4 _0197_
rlabel metal1 s 12972 22202 12972 22202 4 _0198_
rlabel metal1 s 13064 22746 13064 22746 4 _0199_
rlabel metal1 s 10534 22644 10534 22644 4 _0200_
rlabel metal2 s 12282 21250 12282 21250 4 _0201_
rlabel metal1 s 12466 21455 12466 21455 4 _0202_
rlabel metal2 s 13110 21148 13110 21148 4 _0203_
rlabel metal1 s 13984 14926 13984 14926 4 _0204_
rlabel metal2 s 12650 15538 12650 15538 4 _0205_
rlabel metal1 s 13892 15130 13892 15130 4 _0206_
rlabel metal2 s 12834 14076 12834 14076 4 _0207_
rlabel metal1 s 13570 13158 13570 13158 4 _0208_
rlabel metal2 s 13294 12444 13294 12444 4 _0209_
rlabel metal1 s 13018 16014 13018 16014 4 _0210_
rlabel metal1 s 20562 21590 20562 21590 4 _0211_
rlabel metal2 s 10074 20774 10074 20774 4 _0212_
rlabel metal1 s 9890 21012 9890 21012 4 _0213_
rlabel metal2 s 10718 21216 10718 21216 4 _0214_
rlabel metal2 s 9430 21335 9430 21335 4 _0215_
rlabel metal1 s 10902 21522 10902 21522 4 _0216_
rlabel metal1 s 10764 21998 10764 21998 4 _0217_
rlabel metal2 s 12834 22542 12834 22542 4 _0218_
rlabel metal1 s 12834 22474 12834 22474 4 _0219_
rlabel metal1 s 12926 22406 12926 22406 4 _0220_
rlabel metal1 s 13563 21454 13563 21454 4 _0221_
rlabel metal1 s 13432 16014 13432 16014 4 _0222_
rlabel metal1 s 14030 15504 14030 15504 4 _0223_
rlabel metal1 s 13616 15538 13616 15538 4 _0224_
rlabel metal2 s 12926 14382 12926 14382 4 _0225_
rlabel metal2 s 13846 12954 13846 12954 4 _0226_
rlabel metal1 s 14030 12954 14030 12954 4 _0227_
rlabel metal1 s 13984 12614 13984 12614 4 _0228_
rlabel metal2 s 6762 19788 6762 19788 4 _0229_
rlabel metal1 s 8234 19210 8234 19210 4 _0230_
rlabel metal1 s 10718 19890 10718 19890 4 _0231_
rlabel metal2 s 11086 20570 11086 20570 4 _0232_
rlabel metal1 s 12052 18734 12052 18734 4 _0233_
rlabel metal1 s 11730 19346 11730 19346 4 _0234_
rlabel metal2 s 12650 18496 12650 18496 4 _0235_
rlabel metal1 s 13018 19312 13018 19312 4 _0236_
rlabel metal1 s 13279 18802 13279 18802 4 _0237_
rlabel metal1 s 13800 18054 13800 18054 4 _0238_
rlabel metal2 s 13202 18530 13202 18530 4 _0239_
rlabel metal2 s 13938 15028 13938 15028 4 _0240_
rlabel metal2 s 13754 15844 13754 15844 4 _0241_
rlabel metal1 s 13616 17170 13616 17170 4 _0242_
rlabel metal2 s 14122 13906 14122 13906 4 _0243_
rlabel metal2 s 9614 17510 9614 17510 4 _0244_
rlabel metal2 s 9522 18156 9522 18156 4 _0245_
rlabel metal1 s 10810 17850 10810 17850 4 _0246_
rlabel metal1 s 10994 18258 10994 18258 4 _0247_
rlabel metal1 s 12374 18258 12374 18258 4 _0248_
rlabel metal1 s 13018 17510 13018 17510 4 _0249_
rlabel metal1 s 13386 18190 13386 18190 4 _0250_
rlabel metal1 s 12788 17714 12788 17714 4 _0251_
rlabel metal1 s 13892 17714 13892 17714 4 _0252_
rlabel metal1 s 13662 17612 13662 17612 4 _0253_
rlabel metal1 s 15364 12818 15364 12818 4 _0254_
rlabel metal1 s 3956 16762 3956 16762 4 _0255_
rlabel metal1 s 6026 16082 6026 16082 4 _0256_
rlabel metal2 s 7498 16796 7498 16796 4 _0257_
rlabel metal1 s 6670 16082 6670 16082 4 _0258_
rlabel metal1 s 9338 15980 9338 15980 4 _0259_
rlabel metal1 s 8648 16082 8648 16082 4 _0260_
rlabel metal1 s 10442 16218 10442 16218 4 _0261_
rlabel metal1 s 10534 16592 10534 16592 4 _0262_
rlabel metal1 s 12006 16558 12006 16558 4 _0263_
rlabel metal2 s 12190 17340 12190 17340 4 _0264_
rlabel metal2 s 16790 16626 16790 16626 4 _0265_
rlabel metal2 s 16882 16490 16882 16490 4 _0266_
rlabel metal1 s 15364 15538 15364 15538 4 _0267_
rlabel metal2 s 14030 17102 14030 17102 4 _0268_
rlabel metal2 s 15226 16116 15226 16116 4 _0269_
rlabel metal1 s 15042 15470 15042 15470 4 _0270_
rlabel metal1 s 16008 14994 16008 14994 4 _0271_
rlabel metal2 s 15962 14926 15962 14926 4 _0272_
rlabel metal2 s 14766 20638 14766 20638 4 _0273_
rlabel metal1 s 4646 19890 4646 19890 4 _0274_
rlabel metal1 s 5106 19958 5106 19958 4 _0275_
rlabel metal2 s 4922 19006 4922 19006 4 _0276_
rlabel metal2 s 6026 19482 6026 19482 4 _0277_
rlabel metal1 s 5566 19482 5566 19482 4 _0278_
rlabel metal1 s 14674 18836 14674 18836 4 _0279_
rlabel metal2 s 14582 18020 14582 18020 4 _0280_
rlabel metal1 s 16330 18122 16330 18122 4 _0281_
rlabel metal1 s 15824 18258 15824 18258 4 _0282_
rlabel metal2 s 15686 17612 15686 17612 4 _0283_
rlabel metal2 s 15134 16796 15134 16796 4 _0284_
rlabel metal2 s 16054 16524 16054 16524 4 _0285_
rlabel metal2 s 15870 16388 15870 16388 4 _0286_
rlabel metal2 s 16514 16218 16514 16218 4 _0287_
rlabel metal1 s 16438 15946 16438 15946 4 _0288_
rlabel metal2 s 16514 14756 16514 14756 4 _0289_
rlabel metal2 s 16422 14620 16422 14620 4 _0290_
rlabel metal1 s 15410 20944 15410 20944 4 _0291_
rlabel metal2 s 15594 21148 15594 21148 4 _0292_
rlabel metal1 s 15778 21012 15778 21012 4 _0293_
rlabel metal1 s 16928 21658 16928 21658 4 _0294_
rlabel metal1 s 16422 20944 16422 20944 4 _0295_
rlabel metal1 s 16146 19278 16146 19278 4 _0296_
rlabel metal1 s 15962 19414 15962 19414 4 _0297_
rlabel metal1 s 17112 19210 17112 19210 4 _0298_
rlabel metal2 s 16422 18938 16422 18938 4 _0299_
rlabel metal1 s 17296 19482 17296 19482 4 _0300_
rlabel metal1 s 17066 18802 17066 18802 4 _0301_
rlabel metal1 s 16974 18190 16974 18190 4 _0302_
rlabel metal1 s 18492 18802 18492 18802 4 _0303_
rlabel metal2 s 17710 17884 17710 17884 4 _0304_
rlabel metal2 s 17894 17306 17894 17306 4 _0305_
rlabel metal2 s 13202 14620 13202 14620 4 _0306_
rlabel metal1 s 14950 16150 14950 16150 4 _0307_
rlabel metal1 s 17158 15946 17158 15946 4 _0308_
rlabel metal1 s 17066 16184 17066 16184 4 _0309_
rlabel metal1 s 17158 16558 17158 16558 4 _0310_
rlabel metal1 s 18400 16626 18400 16626 4 _0311_
rlabel metal1 s 18814 16762 18814 16762 4 _0312_
rlabel metal1 s 18124 16218 18124 16218 4 _0313_
rlabel metal2 s 18446 15572 18446 15572 4 _0314_
rlabel metal1 s 17304 21318 17304 21318 4 _0315_
rlabel metal2 s 17894 21114 17894 21114 4 _0316_
rlabel metal1 s 17710 21352 17710 21352 4 _0317_
rlabel metal2 s 18078 21114 18078 21114 4 _0318_
rlabel metal2 s 18170 21658 18170 21658 4 _0319_
rlabel metal1 s 17680 19210 17680 19210 4 _0320_
rlabel metal2 s 18078 18972 18078 18972 4 _0321_
rlabel metal1 s 18262 18768 18262 18768 4 _0322_
rlabel metal2 s 18446 17884 18446 17884 4 _0323_
rlabel metal1 s 18860 16014 18860 16014 4 _0324_
rlabel metal2 s 18722 16490 18722 16490 4 _0325_
rlabel metal2 s 20654 22338 20654 22338 4 _0326_
rlabel metal1 s 21758 22610 21758 22610 4 _0327_
rlabel metal1 s 21896 22066 21896 22066 4 _0328_
rlabel metal1 s 20838 21930 20838 21930 4 _0329_
rlabel metal1 s 21114 21998 21114 21998 4 _0330_
rlabel metal1 s 20884 21998 20884 21998 4 _0331_
rlabel metal1 s 20317 21454 20317 21454 4 _0332_
rlabel metal1 s 19550 21522 19550 21522 4 _0333_
rlabel metal2 s 19458 20842 19458 20842 4 _0334_
rlabel metal2 s 19642 20570 19642 20570 4 _0335_
rlabel metal2 s 19182 20060 19182 20060 4 _0336_
rlabel metal1 s 18492 19142 18492 19142 4 _0337_
rlabel metal2 s 18446 19074 18446 19074 4 _0338_
rlabel metal2 s 18722 19584 18722 19584 4 _0339_
rlabel metal1 s 19550 19244 19550 19244 4 _0340_
rlabel metal2 s 19458 19516 19458 19516 4 _0341_
rlabel metal2 s 19734 18836 19734 18836 4 _0342_
rlabel metal1 s 22218 21964 22218 21964 4 _0343_
rlabel metal2 s 22310 21828 22310 21828 4 _0344_
rlabel metal2 s 21758 21182 21758 21182 4 _0345_
rlabel metal2 s 22126 21352 22126 21352 4 _0346_
rlabel metal2 s 21566 20298 21566 20298 4 _0347_
rlabel metal1 s 20976 20570 20976 20570 4 _0348_
rlabel metal1 s 21298 20298 21298 20298 4 _0349_
rlabel metal1 s 20286 17102 20286 17102 4 _0350_
rlabel metal2 s 21298 20400 21298 20400 4 _0351_
rlabel metal2 s 20562 19482 20562 19482 4 _0352_
rlabel metal1 s 21068 18938 21068 18938 4 _0353_
rlabel metal2 s 21298 6188 21298 6188 4 _0354_
rlabel metal1 s 22507 13430 22507 13430 4 _0355_
rlabel metal1 s 22402 13328 22402 13328 4 _0356_
rlabel metal1 s 22080 13362 22080 13362 4 _0357_
rlabel metal1 s 21252 6970 21252 6970 4 _0358_
rlabel metal1 s 21390 8058 21390 8058 4 _0359_
rlabel metal2 s 21758 13124 21758 13124 4 _0360_
rlabel metal2 s 22494 14620 22494 14620 4 _0361_
rlabel metal2 s 21482 14450 21482 14450 4 _0362_
rlabel metal1 s 22080 13974 22080 13974 4 _0363_
rlabel metal1 s 20746 14246 20746 14246 4 _0364_
rlabel metal1 s 20608 13838 20608 13838 4 _0365_
rlabel metal2 s 20194 14144 20194 14144 4 _0366_
rlabel metal1 s 19780 14450 19780 14450 4 _0367_
rlabel metal2 s 19642 14076 19642 14076 4 _0368_
rlabel metal1 s 20102 13906 20102 13906 4 _0369_
rlabel metal1 s 18630 13906 18630 13906 4 _0370_
rlabel metal1 s 18170 12410 18170 12410 4 _0371_
rlabel metal1 s 17580 12614 17580 12614 4 _0372_
rlabel metal1 s 18400 12614 18400 12614 4 _0373_
rlabel metal1 s 18676 12274 18676 12274 4 _0374_
rlabel metal1 s 18308 12954 18308 12954 4 _0375_
rlabel metal2 s 17158 12070 17158 12070 4 _0376_
rlabel metal1 s 17526 11696 17526 11696 4 _0377_
rlabel metal2 s 17342 11866 17342 11866 4 _0378_
rlabel metal1 s 17894 11866 17894 11866 4 _0379_
rlabel metal2 s 15962 10506 15962 10506 4 _0380_
rlabel metal1 s 17066 10132 17066 10132 4 _0381_
rlabel metal1 s 15594 9452 15594 9452 4 _0382_
rlabel metal1 s 16790 9928 16790 9928 4 _0383_
rlabel metal2 s 16882 9826 16882 9826 4 _0384_
rlabel metal2 s 14490 7820 14490 7820 4 _0385_
rlabel metal2 s 14306 7718 14306 7718 4 _0386_
rlabel metal1 s 13754 7956 13754 7956 4 _0387_
rlabel metal2 s 13662 7548 13662 7548 4 _0388_
rlabel metal2 s 14030 7616 14030 7616 4 _0389_
rlabel metal1 s 12374 8432 12374 8432 4 _0390_
rlabel metal2 s 12834 7820 12834 7820 4 _0391_
rlabel metal2 s 13294 7684 13294 7684 4 _0392_
rlabel metal2 s 11086 7242 11086 7242 4 _0393_
rlabel metal1 s 11730 6698 11730 6698 4 _0394_
rlabel metal2 s 11638 8092 11638 8092 4 _0395_
rlabel metal1 s 11224 7378 11224 7378 4 _0396_
rlabel metal1 s 11362 7174 11362 7174 4 _0397_
rlabel metal1 s 9246 7786 9246 7786 4 _0398_
rlabel metal1 s 10580 6698 10580 6698 4 _0399_
rlabel metal2 s 8234 7293 8234 7293 4 _0400_
rlabel metal2 s 8418 7718 8418 7718 4 _0401_
rlabel metal2 s 7958 7616 7958 7616 4 _0402_
rlabel metal2 s 6946 7548 6946 7548 4 _0403_
rlabel metal2 s 7406 7684 7406 7684 4 _0404_
rlabel metal2 s 6302 8874 6302 8874 4 _0405_
rlabel metal1 s 6164 7922 6164 7922 4 _0406_
rlabel metal2 s 6118 8126 6118 8126 4 _0407_
rlabel metal1 s 4922 9962 4922 9962 4 _0408_
rlabel metal2 s 5014 8806 5014 8806 4 _0409_
rlabel metal2 s 5106 9214 5106 9214 4 _0410_
rlabel metal1 s 3910 9894 3910 9894 4 _0411_
rlabel metal1 s 4370 8908 4370 8908 4 _0412_
rlabel metal2 s 5658 4420 5658 4420 4 _0413_
rlabel metal1 s 3220 3706 3220 3706 4 _0414_
rlabel metal1 s 3266 5270 3266 5270 4 _0415_
rlabel metal1 s 4002 8602 4002 8602 4 _0416_
rlabel metal1 s 3941 8364 3941 8364 4 _0417_
rlabel metal1 s 4094 8296 4094 8296 4 _0418_
rlabel metal2 s 5934 8364 5934 8364 4 _0419_
rlabel metal1 s 6601 8058 6601 8058 4 _0420_
rlabel metal1 s 11454 6834 11454 6834 4 _0421_
rlabel metal2 s 13938 7310 13938 7310 4 _0422_
rlabel metal1 s 15548 7718 15548 7718 4 _0423_
rlabel metal1 s 17618 10234 17618 10234 4 _0424_
rlabel metal1 s 19320 12954 19320 12954 4 _0425_
rlabel metal1 s 21666 13906 21666 13906 4 _0426_
rlabel metal1 s 22310 13906 22310 13906 4 _0427_
rlabel metal1 s 21988 13158 21988 13158 4 _0428_
rlabel metal2 s 22034 16966 22034 16966 4 _0429_
rlabel metal2 s 22034 11662 22034 11662 4 _0430_
rlabel metal2 s 4738 4216 4738 4216 4 _0431_
rlabel metal2 s 3450 4080 3450 4080 4 _0432_
rlabel metal2 s 3266 4556 3266 4556 4 _0433_
rlabel metal2 s 2346 7174 2346 7174 4 _0434_
rlabel metal1 s 2384 6970 2384 6970 4 _0435_
rlabel metal1 s 2944 6834 2944 6834 4 _0436_
rlabel metal2 s 2990 7174 2990 7174 4 _0437_
rlabel metal1 s 4784 5814 4784 5814 4 _0438_
rlabel metal1 s 4692 6426 4692 6426 4 _0439_
rlabel metal1 s 5934 6426 5934 6426 4 _0440_
rlabel metal1 s 5704 5882 5704 5882 4 _0441_
rlabel metal1 s 6716 6222 6716 6222 4 _0442_
rlabel metal1 s 6716 6426 6716 6426 4 _0443_
rlabel metal1 s 10166 5814 10166 5814 4 _0444_
rlabel metal2 s 8050 5712 8050 5712 4 _0445_
rlabel metal2 s 8786 5440 8786 5440 4 _0446_
rlabel metal1 s 8940 5066 8940 5066 4 _0447_
rlabel metal1 s 10488 4522 10488 4522 4 _0448_
rlabel metal2 s 10350 4998 10350 4998 4 _0449_
rlabel metal1 s 11592 5678 11592 5678 4 _0450_
rlabel metal1 s 11684 4114 11684 4114 4 _0451_
rlabel metal2 s 12742 5440 12742 5440 4 _0452_
rlabel metal1 s 12896 5066 12896 5066 4 _0453_
rlabel metal1 s 14122 6086 14122 6086 4 _0454_
rlabel metal1 s 13892 5542 13892 5542 4 _0455_
rlabel metal2 s 16874 8058 16874 8058 4 _0456_
rlabel metal2 s 15226 5814 15226 5814 4 _0457_
rlabel metal2 s 16238 6800 16238 6800 4 _0458_
rlabel metal1 s 16200 6154 16200 6154 4 _0459_
rlabel metal1 s 15134 8364 15134 8364 4 _0460_
rlabel metal1 s 15824 8058 15824 8058 4 _0461_
rlabel metal2 s 18078 10710 18078 10710 4 _0462_
rlabel metal1 s 16698 9146 16698 9146 4 _0463_
rlabel metal1 s 18906 9622 18906 9622 4 _0464_
rlabel metal1 s 19212 9418 19212 9418 4 _0465_
rlabel metal1 s 20470 11186 20470 11186 4 _0466_
rlabel metal2 s 18538 10506 18538 10506 4 _0467_
rlabel metal2 s 19550 10268 19550 10268 4 _0468_
rlabel metal2 s 19918 10438 19918 10438 4 _0469_
rlabel metal2 s 19550 11968 19550 11968 4 _0470_
rlabel metal1 s 20240 11866 20240 11866 4 _0471_
rlabel metal1 s 20792 9486 20792 9486 4 _0472_
rlabel metal1 s 21344 10982 21344 10982 4 _0473_
rlabel metal1 s 21344 9962 21344 9962 4 _0474_
rlabel metal1 s 21344 9690 21344 9690 4 _0475_
rlabel metal1 s 21896 8534 21896 8534 4 _0476_
rlabel metal2 s 22034 9282 22034 9282 4 _0477_
rlabel metal1 s 22218 5848 22218 5848 4 _0478_
rlabel metal2 s 21390 7616 21390 7616 4 _0479_
rlabel metal2 s 22586 6052 22586 6052 4 _0480_
rlabel metal1 s 20700 6290 20700 6290 4 _0481_
rlabel metal1 s 20470 5066 20470 5066 4 _0482_
rlabel metal1 s 19550 5066 19550 5066 4 _0483_
rlabel metal2 s 19826 6868 19826 6868 4 _0484_
rlabel metal1 s 19136 6154 19136 6154 4 _0485_
rlabel metal1 s 19642 7344 19642 7344 4 _0486_
rlabel metal1 s 19136 7514 19136 7514 4 _0487_
rlabel metal1 s 18706 7242 18706 7242 4 _0488_
rlabel metal1 s 21804 16218 21804 16218 4 _0489_
rlabel metal2 s 23046 3961 23046 3961 4 clk_in
rlabel metal2 s 23046 19465 23046 19465 4 clk_out
rlabel metal1 s 2714 4250 2714 4250 4 count\[0\]
rlabel metal2 s 10074 4216 10074 4216 4 count\[10\]
rlabel metal1 s 10580 5746 10580 5746 4 count\[11\]
rlabel metal1 s 11224 5882 11224 5882 4 count\[12\]
rlabel metal2 s 13018 6528 13018 6528 4 count\[13\]
rlabel metal2 s 14306 5372 14306 5372 4 count\[14\]
rlabel metal2 s 14950 5746 14950 5746 4 count\[15\]
rlabel metal2 s 15870 9758 15870 9758 4 count\[16\]
rlabel metal2 s 16606 9792 16606 9792 4 count\[17\]
rlabel metal1 s 16698 12376 16698 12376 4 count\[18\]
rlabel metal1 s 17526 12716 17526 12716 4 count\[19\]
rlabel metal1 s 3542 4012 3542 4012 4 count\[1\]
rlabel metal2 s 18446 11628 18446 11628 4 count\[20\]
rlabel metal1 s 19458 13838 19458 13838 4 count\[21\]
rlabel metal2 s 21114 14178 21114 14178 4 count\[22\]
rlabel metal2 s 21574 13129 21574 13129 4 count\[23\]
rlabel metal2 s 22218 12920 22218 12920 4 count\[24\]
rlabel metal1 s 22402 13804 22402 13804 4 count\[25\]
rlabel metal1 s 21666 7956 21666 7956 4 count\[26\]
rlabel metal1 s 22402 5712 22402 5712 4 count\[27\]
rlabel metal2 s 20930 4964 20930 4964 4 count\[28\]
rlabel metal1 s 20194 6698 20194 6698 4 count\[29\]
rlabel metal1 s 3312 4046 3312 4046 4 count\[2\]
rlabel metal1 s 20102 6868 20102 6868 4 count\[30\]
rlabel metal1 s 20838 7786 20838 7786 4 count\[31\]
rlabel metal1 s 4002 4794 4002 4794 4 count\[3\]
rlabel metal2 s 3358 7174 3358 7174 4 count\[4\]
rlabel metal1 s 3358 6630 3358 6630 4 count\[5\]
rlabel metal1 s 4692 8330 4692 8330 4 count\[6\]
rlabel metal1 s 5934 6222 5934 6222 4 count\[7\]
rlabel metal1 s 7176 6222 7176 6222 4 count\[8\]
rlabel metal1 s 7636 5882 7636 5882 4 count\[9\]
rlabel metal2 s 22862 4352 22862 4352 4 net1
rlabel metal1 s 22770 22168 22770 22168 4 net10
rlabel metal1 s 2760 5338 2760 5338 4 net11
rlabel metal1 s 20286 12308 20286 12308 4 net12
rlabel metal1 s 13110 5814 13110 5814 4 net13
rlabel metal1 s 22172 11050 22172 11050 4 net14
rlabel metal1 s 13524 12818 13524 12818 4 net15
rlabel metal1 s 5842 11118 5842 11118 4 net16
rlabel metal1 s 14858 21862 14858 21862 4 net17
rlabel metal1 s 4002 23188 4002 23188 4 net18
rlabel metal2 s 2898 14144 2898 14144 4 net19
rlabel metal1 s 22770 17000 22770 17000 4 net2
rlabel metal1 s 3542 22984 3542 22984 4 net20
rlabel metal1 s 15548 14450 15548 14450 4 net21
rlabel metal2 s 3266 11900 3266 11900 4 net22
rlabel metal1 s 2668 4658 2668 4658 4 net23
rlabel metal1 s 6394 4590 6394 4590 4 net24
rlabel metal1 s 4738 11730 4738 11730 4 net25
rlabel metal1 s 19642 10574 19642 10574 4 net26
rlabel metal1 s 20700 6154 20700 6154 4 net27
rlabel metal2 s 22310 18938 22310 18938 4 net28
rlabel metal2 s 22678 17714 22678 17714 4 net29
rlabel metal2 s 3082 22746 3082 22746 4 net3
rlabel metal1 s 3404 23222 3404 23222 4 net4
rlabel metal1 s 5152 23154 5152 23154 4 net5
rlabel metal2 s 4738 22644 4738 22644 4 net6
rlabel metal1 s 16882 21454 16882 21454 4 net7
rlabel metal1 s 22310 22066 22310 22066 4 net8
rlabel metal1 s 21896 21454 21896 21454 4 net9
rlabel metal2 s 23046 12019 23046 12019 4 nrst
rlabel metal2 s 1794 23443 1794 23443 4 scale[0]
rlabel metal1 s 5382 23188 5382 23188 4 scale[1]
rlabel metal1 s 7728 23154 7728 23154 4 scale[2]
rlabel metal1 s 10810 23222 10810 23222 4 scale[3]
rlabel metal2 s 13570 23443 13570 23443 4 scale[4]
rlabel metal2 s 16514 23443 16514 23443 4 scale[5]
rlabel metal2 s 19458 23443 19458 23443 4 scale[6]
rlabel metal1 s 22356 23154 22356 23154 4 scale[7]
rlabel metal1 s 22586 17102 22586 17102 4 signal_clk_out
rlabel metal1 s 7636 10234 7636 10234 4 true_scale\[10\]
rlabel metal2 s 8786 9248 8786 9248 4 true_scale\[11\]
rlabel metal2 s 10810 9248 10810 9248 4 true_scale\[12\]
rlabel metal1 s 10764 10778 10764 10778 4 true_scale\[13\]
rlabel metal2 s 11270 10982 11270 10982 4 true_scale\[14\]
rlabel metal1 s 13800 11118 13800 11118 4 true_scale\[15\]
rlabel metal1 s 12903 9690 12903 9690 4 true_scale\[16\]
rlabel metal1 s 13386 9520 13386 9520 4 true_scale\[17\]
rlabel metal1 s 15640 12682 15640 12682 4 true_scale\[18\]
rlabel metal1 s 16192 14042 16192 14042 4 true_scale\[19\]
rlabel metal2 s 17526 13906 17526 13906 4 true_scale\[20\]
rlabel metal2 s 19458 14892 19458 14892 4 true_scale\[21\]
rlabel metal1 s 19090 15946 19090 15946 4 true_scale\[22\]
rlabel metal1 s 20378 14858 20378 14858 4 true_scale\[23\]
rlabel metal1 s 20884 16966 20884 16966 4 true_scale\[24\]
rlabel metal2 s 22310 15742 22310 15742 4 true_scale\[25\]
rlabel metal1 s 21206 18598 21206 18598 4 true_scale\[26\]
rlabel metal1 s 3312 11866 3312 11866 4 true_scale\[5\]
rlabel metal1 s 3496 10030 3496 10030 4 true_scale\[6\]
rlabel metal1 s 4876 11322 4876 11322 4 true_scale\[7\]
rlabel metal1 s 4646 9554 4646 9554 4 true_scale\[8\]
rlabel metal2 s 6762 10982 6762 10982 4 true_scale\[9\]
flabel metal4 s 4316 496 4636 23440 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 3656 496 3976 23440 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 23600 3816 24000 3936 0 FreeSans 600 0 0 0 clk_in
port 3 nsew
flabel metal3 s 23600 19592 24000 19712 0 FreeSans 600 0 0 0 clk_out
port 4 nsew
flabel metal3 s 23600 11704 24000 11824 0 FreeSans 600 0 0 0 nrst
port 5 nsew
flabel metal2 s 1674 23600 1730 24000 0 FreeSans 280 90 0 0 scale[0]
port 6 nsew
flabel metal2 s 4618 23600 4674 24000 0 FreeSans 280 90 0 0 scale[1]
port 7 nsew
flabel metal2 s 7562 23600 7618 24000 0 FreeSans 280 90 0 0 scale[2]
port 8 nsew
flabel metal2 s 10506 23600 10562 24000 0 FreeSans 280 90 0 0 scale[3]
port 9 nsew
flabel metal2 s 13450 23600 13506 24000 0 FreeSans 280 90 0 0 scale[4]
port 10 nsew
flabel metal2 s 16394 23600 16450 24000 0 FreeSans 280 90 0 0 scale[5]
port 11 nsew
flabel metal2 s 19338 23600 19394 24000 0 FreeSans 280 90 0 0 scale[6]
port 12 nsew
flabel metal2 s 22282 23600 22338 24000 0 FreeSans 280 90 0 0 scale[7]
port 13 nsew
<< properties >>
string FIXED_BBOX 0 0 24000 24000
string GDS_END 1764632
string GDS_FILE clock_divider.gds
string GDS_START 501286
<< end >>
