magic
tech sky130A
timestamp 1701394307
<< pwell >>
rect -848 -855 848 855
<< nmos >>
rect -750 -750 750 750
<< ndiff >>
rect -779 744 -750 750
rect -779 -744 -773 744
rect -756 -744 -750 744
rect -779 -750 -750 -744
rect 750 744 779 750
rect 750 -744 756 744
rect 773 -744 779 744
rect 750 -750 779 -744
<< ndiffc >>
rect -773 -744 -756 744
rect 756 -744 773 744
<< psubdiff >>
rect -830 820 -782 837
rect 782 820 830 837
rect -830 789 -813 820
rect 813 789 830 820
rect -830 -820 -813 -789
rect 813 -820 830 -789
rect -830 -837 -782 -820
rect 782 -837 830 -820
<< psubdiffcont >>
rect -782 820 782 837
rect -830 -789 -813 789
rect 813 -789 830 789
rect -782 -837 782 -820
<< poly >>
rect -750 786 750 794
rect -750 769 -742 786
rect 742 769 750 786
rect -750 750 750 769
rect -750 -769 750 -750
rect -750 -786 -742 -769
rect 742 -786 750 -769
rect -750 -794 750 -786
<< polycont >>
rect -742 769 742 786
rect -742 -786 742 -769
<< locali >>
rect -830 820 -782 837
rect 782 820 830 837
rect -830 789 -813 820
rect 813 789 830 820
rect -750 769 -742 786
rect 742 769 750 786
rect -773 744 -756 752
rect -773 -752 -756 -744
rect 756 744 773 752
rect 756 -752 773 -744
rect -750 -786 -742 -769
rect 742 -786 750 -769
rect -830 -820 -813 -789
rect 813 -820 830 -789
rect -830 -837 -782 -820
rect 782 -837 830 -820
<< viali >>
rect -742 769 742 786
rect -773 -744 -756 744
rect 756 -744 773 744
rect -742 -786 742 -769
<< metal1 >>
rect -748 786 748 789
rect -748 769 -742 786
rect 742 769 748 786
rect -748 766 748 769
rect -776 744 -753 750
rect -776 -744 -773 744
rect -756 -744 -753 744
rect -776 -750 -753 -744
rect 753 744 776 750
rect 753 -744 756 744
rect 773 -744 776 744
rect 753 -750 776 -744
rect -748 -769 748 -766
rect -748 -786 -742 -769
rect 742 -786 748 -769
rect -748 -789 748 -786
<< properties >>
string FIXED_BBOX -821 -828 821 828
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 15 l 15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
