magic
tech sky130A
magscale 1 2
timestamp 1700708449
<< metal3 >>
rect -3186 1112 3186 1140
rect -3186 -1112 3102 1112
rect 3166 -1112 3186 1112
rect -3186 -1140 3186 -1112
<< via3 >>
rect 3102 -1112 3166 1112
<< mimcap >>
rect -3146 1060 2854 1100
rect -3146 -1060 -3106 1060
rect 2814 -1060 2854 1060
rect -3146 -1100 2854 -1060
<< mimcapcontact >>
rect -3106 -1060 2814 1060
<< metal4 >>
rect 3086 1112 3182 1128
rect -3107 1060 2815 1061
rect -3107 -1060 -3106 1060
rect 2814 -1060 2815 1060
rect -3107 -1061 2815 -1060
rect 3086 -1112 3102 1112
rect 3166 -1112 3182 1112
rect 3086 -1128 3182 -1112
<< properties >>
string FIXED_BBOX -3186 -1140 2894 1140
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30 l 11 val 675.58 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
