magic
tech sky130A
magscale 1 2
timestamp 1700708449
<< metal4 >>
rect -3349 1039 3349 1080
rect -3349 -1039 3093 1039
rect 3329 -1039 3349 1039
rect -3349 -1080 3349 -1039
<< via4 >>
rect 3093 -1039 3329 1039
<< mimcap2 >>
rect -3269 960 2731 1000
rect -3269 -960 -3229 960
rect 2691 -960 2731 960
rect -3269 -1000 2731 -960
<< mimcap2contact >>
rect -3229 -960 2691 960
<< metal5 >>
rect 3051 1039 3371 1081
rect -3253 960 2715 984
rect -3253 -960 -3229 960
rect 2691 -960 2715 960
rect -3253 -984 2715 -960
rect 3051 -1039 3093 1039
rect 3329 -1039 3371 1039
rect 3051 -1081 3371 -1039
<< properties >>
string FIXED_BBOX -3349 -1080 2811 1080
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 30 l 10 val 615.2 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
