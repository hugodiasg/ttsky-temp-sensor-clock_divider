magic
tech sky130A
magscale 1 2
timestamp 1700747326
<< pwell >>
rect -1596 -1210 1596 1210
<< nmos >>
rect -1400 -1000 1400 1000
<< ndiff >>
rect -1458 988 -1400 1000
rect -1458 -988 -1446 988
rect -1412 -988 -1400 988
rect -1458 -1000 -1400 -988
rect 1400 988 1458 1000
rect 1400 -988 1412 988
rect 1446 -988 1458 988
rect 1400 -1000 1458 -988
<< ndiffc >>
rect -1446 -988 -1412 988
rect 1412 -988 1446 988
<< psubdiff >>
rect -1560 1140 -1464 1174
rect 1464 1140 1560 1174
rect -1560 1078 -1526 1140
rect 1526 1078 1560 1140
rect -1560 -1140 -1526 -1078
rect 1526 -1140 1560 -1078
rect -1560 -1174 -1464 -1140
rect 1464 -1174 1560 -1140
<< psubdiffcont >>
rect -1464 1140 1464 1174
rect -1560 -1078 -1526 1078
rect 1526 -1078 1560 1078
rect -1464 -1174 1464 -1140
<< poly >>
rect -1400 1072 1400 1088
rect -1400 1038 -1384 1072
rect 1384 1038 1400 1072
rect -1400 1000 1400 1038
rect -1400 -1038 1400 -1000
rect -1400 -1072 -1384 -1038
rect 1384 -1072 1400 -1038
rect -1400 -1088 1400 -1072
<< polycont >>
rect -1384 1038 1384 1072
rect -1384 -1072 1384 -1038
<< locali >>
rect -1560 1140 -1464 1174
rect 1464 1140 1560 1174
rect -1560 1078 -1526 1140
rect 1526 1078 1560 1140
rect -1400 1038 -1384 1072
rect 1384 1038 1400 1072
rect -1446 988 -1412 1004
rect -1446 -1004 -1412 -988
rect 1412 988 1446 1004
rect 1412 -1004 1446 -988
rect -1400 -1072 -1384 -1038
rect 1384 -1072 1400 -1038
rect -1560 -1140 -1526 -1078
rect 1526 -1140 1560 -1078
rect -1560 -1174 -1464 -1140
rect 1464 -1174 1560 -1140
<< viali >>
rect -1384 1038 1384 1072
rect -1446 -971 -1412 17
rect 1412 -17 1446 971
rect -1384 -1072 1384 -1038
<< metal1 >>
rect -1396 1072 1396 1078
rect -1396 1038 -1384 1072
rect 1384 1038 1396 1072
rect -1396 1032 1396 1038
rect 1406 971 1452 983
rect -1452 17 -1406 29
rect -1452 -971 -1446 17
rect -1412 -971 -1406 17
rect 1406 -17 1412 971
rect 1446 -17 1452 971
rect 1406 -29 1452 -17
rect -1452 -983 -1406 -971
rect -1396 -1038 1396 -1032
rect -1396 -1072 -1384 -1038
rect 1384 -1072 1396 -1038
rect -1396 -1078 1396 -1072
<< properties >>
string FIXED_BBOX -1543 -1157 1543 1157
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 10 l 14 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc -50 viadrn +50 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
