magic
tech sky130A
magscale 1 2
timestamp 1700703435
<< metal4 >>
rect -2349 2239 2349 2280
rect -2349 -2239 2093 2239
rect 2329 -2239 2349 2239
rect -2349 -2280 2349 -2239
<< via4 >>
rect 2093 -2239 2329 2239
<< mimcap2 >>
rect -2269 2160 1731 2200
rect -2269 -2160 -2229 2160
rect 1691 -2160 1731 2160
rect -2269 -2200 1731 -2160
<< mimcap2contact >>
rect -2229 -2160 1691 2160
<< metal5 >>
rect 2051 2239 2371 2281
rect -2253 2160 1715 2184
rect -2253 -2160 -2229 2160
rect 1691 -2160 1715 2160
rect -2253 -2184 1715 -2160
rect 2051 -2239 2093 2239
rect 2329 -2239 2371 2239
rect 2051 -2281 2371 -2239
<< properties >>
string FIXED_BBOX -2349 -2280 1811 2280
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 20 l 22 val 895.96 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
