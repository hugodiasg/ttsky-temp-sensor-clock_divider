magic
tech sky130A
timestamp 1699933188
<< pwell >>
rect -898 -455 898 455
<< nmos >>
rect -800 -350 800 350
<< ndiff >>
rect -829 344 -800 350
rect -829 -344 -823 344
rect -806 -344 -800 344
rect -829 -350 -800 -344
rect 800 344 829 350
rect 800 -344 806 344
rect 823 -344 829 344
rect 800 -350 829 -344
<< ndiffc >>
rect -823 -344 -806 344
rect 806 -344 823 344
<< psubdiff >>
rect -880 420 -832 437
rect 832 420 880 437
rect -880 389 -863 420
rect 863 389 880 420
rect -880 -420 -863 -389
rect 863 -420 880 -389
rect -880 -437 -832 -420
rect 832 -437 880 -420
<< psubdiffcont >>
rect -832 420 832 437
rect -880 -389 -863 389
rect 863 -389 880 389
rect -832 -437 832 -420
<< poly >>
rect -800 386 800 394
rect -800 369 -792 386
rect 792 369 800 386
rect -800 350 800 369
rect -800 -369 800 -350
rect -800 -386 -792 -369
rect 792 -386 800 -369
rect -800 -394 800 -386
<< polycont >>
rect -792 369 792 386
rect -792 -386 792 -369
<< locali >>
rect -880 420 -832 437
rect 832 420 880 437
rect -880 389 -863 420
rect 863 389 880 420
rect -800 369 -792 386
rect 792 369 800 386
rect -823 344 -806 352
rect -823 -352 -806 -344
rect 806 344 823 352
rect 806 -352 823 -344
rect -800 -386 -792 -369
rect 792 -386 800 -369
rect -880 -420 -863 -389
rect 863 -420 880 -389
rect -880 -437 -832 -420
rect 832 -437 880 -420
<< viali >>
rect -792 369 792 386
rect -823 -344 -806 344
rect 806 -344 823 344
rect -792 -386 792 -369
<< metal1 >>
rect -798 386 798 389
rect -798 369 -792 386
rect 792 369 798 386
rect -798 366 798 369
rect -826 344 -803 350
rect -826 -344 -823 344
rect -806 -344 -803 344
rect -826 -350 -803 -344
rect 803 344 826 350
rect 803 -344 806 344
rect 823 -344 826 344
rect 803 -350 826 -344
rect -798 -369 798 -366
rect -798 -386 -792 -369
rect 792 -386 798 -369
rect -798 -389 798 -386
<< properties >>
string FIXED_BBOX -871 -428 871 428
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 7 l 16 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
