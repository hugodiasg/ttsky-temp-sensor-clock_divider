magic
tech sky130A
magscale 1 2
timestamp 1699932112
<< nwell >>
rect -581 -300 581 300
<< pmos >>
rect -487 -200 -287 200
rect -229 -200 -29 200
rect 29 -200 229 200
rect 287 -200 487 200
<< pdiff >>
rect -545 188 -487 200
rect -545 -188 -533 188
rect -499 -188 -487 188
rect -545 -200 -487 -188
rect -287 188 -229 200
rect -287 -188 -275 188
rect -241 -188 -229 188
rect -287 -200 -229 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 229 188 287 200
rect 229 -188 241 188
rect 275 -188 287 188
rect 229 -200 287 -188
rect 487 188 545 200
rect 487 -188 499 188
rect 533 -188 545 188
rect 487 -200 545 -188
<< pdiffc >>
rect -533 -188 -499 188
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect 499 -188 533 188
<< poly >>
rect -487 281 -287 297
rect -487 247 -471 281
rect -303 247 -287 281
rect -487 200 -287 247
rect -229 281 -29 297
rect -229 247 -213 281
rect -45 247 -29 281
rect -229 200 -29 247
rect 29 281 229 297
rect 29 247 45 281
rect 213 247 229 281
rect 29 200 229 247
rect 287 281 487 297
rect 287 247 303 281
rect 471 247 487 281
rect 287 200 487 247
rect -487 -247 -287 -200
rect -487 -281 -471 -247
rect -303 -281 -287 -247
rect -487 -297 -287 -281
rect -229 -247 -29 -200
rect -229 -281 -213 -247
rect -45 -281 -29 -247
rect -229 -297 -29 -281
rect 29 -247 229 -200
rect 29 -281 45 -247
rect 213 -281 229 -247
rect 29 -297 229 -281
rect 287 -247 487 -200
rect 287 -281 303 -247
rect 471 -281 487 -247
rect 287 -297 487 -281
<< polycont >>
rect -471 247 -303 281
rect -213 247 -45 281
rect 45 247 213 281
rect 303 247 471 281
rect -471 -281 -303 -247
rect -213 -281 -45 -247
rect 45 -281 213 -247
rect 303 -281 471 -247
<< locali >>
rect -487 247 -471 281
rect -303 247 -287 281
rect -229 247 -213 281
rect -45 247 -29 281
rect 29 247 45 281
rect 213 247 229 281
rect 287 247 303 281
rect 471 247 487 281
rect -533 188 -499 204
rect -533 -204 -499 -188
rect -275 188 -241 204
rect -275 -204 -241 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 241 188 275 204
rect 241 -204 275 -188
rect 499 188 533 204
rect 499 -204 533 -188
rect -487 -281 -471 -247
rect -303 -281 -287 -247
rect -229 -281 -213 -247
rect -45 -281 -29 -247
rect 29 -281 45 -247
rect 213 -281 229 -247
rect 287 -281 303 -247
rect 471 -281 487 -247
<< viali >>
rect -471 247 -303 281
rect -213 247 -45 281
rect 45 247 213 281
rect 303 247 471 281
rect -533 -171 -499 17
rect -275 -17 -241 171
rect -17 -171 17 17
rect 241 -17 275 171
rect 499 -171 533 17
rect -471 -281 -303 -247
rect -213 -281 -45 -247
rect 45 -281 213 -247
rect 303 -281 471 -247
<< metal1 >>
rect -483 281 -291 287
rect -483 247 -471 281
rect -303 247 -291 281
rect -483 241 -291 247
rect -225 281 -33 287
rect -225 247 -213 281
rect -45 247 -33 281
rect -225 241 -33 247
rect 33 281 225 287
rect 33 247 45 281
rect 213 247 225 281
rect 33 241 225 247
rect 291 281 483 287
rect 291 247 303 281
rect 471 247 483 281
rect 291 241 483 247
rect -281 171 -235 183
rect -539 17 -493 29
rect -539 -171 -533 17
rect -499 -171 -493 17
rect -281 -17 -275 171
rect -241 -17 -235 171
rect 235 171 281 183
rect -281 -29 -235 -17
rect -23 17 23 29
rect -539 -183 -493 -171
rect -23 -171 -17 17
rect 17 -171 23 17
rect 235 -17 241 171
rect 275 -17 281 171
rect 235 -29 281 -17
rect 493 17 539 29
rect -23 -183 23 -171
rect 493 -171 499 17
rect 533 -171 539 17
rect 493 -183 539 -171
rect -483 -247 -291 -241
rect -483 -281 -471 -247
rect -303 -281 -291 -247
rect -483 -287 -291 -281
rect -225 -247 -33 -241
rect -225 -281 -213 -247
rect -45 -281 -33 -247
rect -225 -287 -33 -281
rect 33 -247 225 -241
rect 33 -281 45 -247
rect 213 -281 225 -247
rect 33 -287 225 -281
rect 291 -247 483 -241
rect 291 -281 303 -247
rect 471 -281 483 -247
rect 291 -287 483 -281
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 1 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc -50 viadrn +50 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
