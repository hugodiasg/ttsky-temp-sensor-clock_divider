magic
tech sky130A
magscale 1 2
timestamp 1700746600
<< nwell >>
rect -968 -200 968 200
<< pmos >>
rect -874 -100 -674 100
rect -616 -100 -416 100
rect -358 -100 -158 100
rect -100 -100 100 100
rect 158 -100 358 100
rect 416 -100 616 100
rect 674 -100 874 100
<< pdiff >>
rect -932 88 -874 100
rect -932 -88 -920 88
rect -886 -88 -874 88
rect -932 -100 -874 -88
rect -674 88 -616 100
rect -674 -88 -662 88
rect -628 -88 -616 88
rect -674 -100 -616 -88
rect -416 88 -358 100
rect -416 -88 -404 88
rect -370 -88 -358 88
rect -416 -100 -358 -88
rect -158 88 -100 100
rect -158 -88 -146 88
rect -112 -88 -100 88
rect -158 -100 -100 -88
rect 100 88 158 100
rect 100 -88 112 88
rect 146 -88 158 88
rect 100 -100 158 -88
rect 358 88 416 100
rect 358 -88 370 88
rect 404 -88 416 88
rect 358 -100 416 -88
rect 616 88 674 100
rect 616 -88 628 88
rect 662 -88 674 88
rect 616 -100 674 -88
rect 874 88 932 100
rect 874 -88 886 88
rect 920 -88 932 88
rect 874 -100 932 -88
<< pdiffc >>
rect -920 -88 -886 88
rect -662 -88 -628 88
rect -404 -88 -370 88
rect -146 -88 -112 88
rect 112 -88 146 88
rect 370 -88 404 88
rect 628 -88 662 88
rect 886 -88 920 88
<< poly >>
rect -874 181 -674 197
rect -874 147 -858 181
rect -690 147 -674 181
rect -874 100 -674 147
rect -616 181 -416 197
rect -616 147 -600 181
rect -432 147 -416 181
rect -616 100 -416 147
rect -358 181 -158 197
rect -358 147 -342 181
rect -174 147 -158 181
rect -358 100 -158 147
rect -100 181 100 197
rect -100 147 -84 181
rect 84 147 100 181
rect -100 100 100 147
rect 158 181 358 197
rect 158 147 174 181
rect 342 147 358 181
rect 158 100 358 147
rect 416 181 616 197
rect 416 147 432 181
rect 600 147 616 181
rect 416 100 616 147
rect 674 181 874 197
rect 674 147 690 181
rect 858 147 874 181
rect 674 100 874 147
rect -874 -147 -674 -100
rect -874 -181 -858 -147
rect -690 -181 -674 -147
rect -874 -197 -674 -181
rect -616 -147 -416 -100
rect -616 -181 -600 -147
rect -432 -181 -416 -147
rect -616 -197 -416 -181
rect -358 -147 -158 -100
rect -358 -181 -342 -147
rect -174 -181 -158 -147
rect -358 -197 -158 -181
rect -100 -147 100 -100
rect -100 -181 -84 -147
rect 84 -181 100 -147
rect -100 -197 100 -181
rect 158 -147 358 -100
rect 158 -181 174 -147
rect 342 -181 358 -147
rect 158 -197 358 -181
rect 416 -147 616 -100
rect 416 -181 432 -147
rect 600 -181 616 -147
rect 416 -197 616 -181
rect 674 -147 874 -100
rect 674 -181 690 -147
rect 858 -181 874 -147
rect 674 -197 874 -181
<< polycont >>
rect -858 147 -690 181
rect -600 147 -432 181
rect -342 147 -174 181
rect -84 147 84 181
rect 174 147 342 181
rect 432 147 600 181
rect 690 147 858 181
rect -858 -181 -690 -147
rect -600 -181 -432 -147
rect -342 -181 -174 -147
rect -84 -181 84 -147
rect 174 -181 342 -147
rect 432 -181 600 -147
rect 690 -181 858 -147
<< locali >>
rect -874 147 -858 181
rect -690 147 -674 181
rect -616 147 -600 181
rect -432 147 -416 181
rect -358 147 -342 181
rect -174 147 -158 181
rect -100 147 -84 181
rect 84 147 100 181
rect 158 147 174 181
rect 342 147 358 181
rect 416 147 432 181
rect 600 147 616 181
rect 674 147 690 181
rect 858 147 874 181
rect -920 88 -886 104
rect -920 -104 -886 -88
rect -662 88 -628 104
rect -662 -104 -628 -88
rect -404 88 -370 104
rect -404 -104 -370 -88
rect -146 88 -112 104
rect -146 -104 -112 -88
rect 112 88 146 104
rect 112 -104 146 -88
rect 370 88 404 104
rect 370 -104 404 -88
rect 628 88 662 104
rect 628 -104 662 -88
rect 886 88 920 104
rect 886 -104 920 -88
rect -874 -181 -858 -147
rect -690 -181 -674 -147
rect -616 -181 -600 -147
rect -432 -181 -416 -147
rect -358 -181 -342 -147
rect -174 -181 -158 -147
rect -100 -181 -84 -147
rect 84 -181 100 -147
rect 158 -181 174 -147
rect 342 -181 358 -147
rect 416 -181 432 -147
rect 600 -181 616 -147
rect 674 -181 690 -147
rect 858 -181 874 -147
<< viali >>
rect -920 -71 -886 17
rect -662 -17 -628 71
rect -404 -71 -370 17
rect -146 -17 -112 71
rect 112 -71 146 17
rect 370 -17 404 71
rect 628 -71 662 17
rect 886 -17 920 71
<< metal1 >>
rect -668 71 -622 83
rect -926 17 -880 29
rect -926 -71 -920 17
rect -886 -71 -880 17
rect -668 -17 -662 71
rect -628 -17 -622 71
rect -152 71 -106 83
rect -668 -29 -622 -17
rect -410 17 -364 29
rect -926 -83 -880 -71
rect -410 -71 -404 17
rect -370 -71 -364 17
rect -152 -17 -146 71
rect -112 -17 -106 71
rect 364 71 410 83
rect -152 -29 -106 -17
rect 106 17 152 29
rect -410 -83 -364 -71
rect 106 -71 112 17
rect 146 -71 152 17
rect 364 -17 370 71
rect 404 -17 410 71
rect 880 71 926 83
rect 364 -29 410 -17
rect 622 17 668 29
rect 106 -83 152 -71
rect 622 -71 628 17
rect 662 -71 668 17
rect 880 -17 886 71
rect 920 -17 926 71
rect 880 -29 926 -17
rect 622 -83 668 -71
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.0 l 1.0 m 1 nf 7 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc -50 viadrn +50 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
