magic
tech sky130A
magscale 1 2
timestamp 1700708449
<< metal4 >>
rect -3349 739 3349 780
rect -3349 -739 3093 739
rect 3329 -739 3349 739
rect -3349 -780 3349 -739
<< via4 >>
rect 3093 -739 3329 739
<< mimcap2 >>
rect -3269 660 2731 700
rect -3269 -660 -3229 660
rect 2691 -660 2731 660
rect -3269 -700 2731 -660
<< mimcap2contact >>
rect -3229 -660 2691 660
<< metal5 >>
rect 3051 739 3371 781
rect -3253 660 2715 684
rect -3253 -660 -3229 660
rect 2691 -660 2715 660
rect -3253 -684 2715 -660
rect 3051 -739 3093 739
rect 3329 -739 3371 739
rect 3051 -781 3371 -739
<< properties >>
string FIXED_BBOX -3349 -780 2811 780
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 30 l 7 val 434.06 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
