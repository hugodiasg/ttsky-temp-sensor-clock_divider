magic
tech sky130A
magscale 1 2
timestamp 1700703435
<< metal4 >>
rect -2049 3039 2049 3080
rect -2049 -3039 1793 3039
rect 2029 -3039 2049 3039
rect -2049 -3080 2049 -3039
<< via4 >>
rect 1793 -3039 2029 3039
<< mimcap2 >>
rect -1969 2960 1431 3000
rect -1969 -2960 -1929 2960
rect 1391 -2960 1431 2960
rect -1969 -3000 1431 -2960
<< mimcap2contact >>
rect -1929 -2960 1391 2960
<< metal5 >>
rect 1751 3039 2071 3081
rect -1953 2960 1415 2984
rect -1953 -2960 -1929 2960
rect 1391 -2960 1415 2960
rect -1953 -2984 1415 -2960
rect 1751 -3039 1793 3039
rect 2029 -3039 2071 3039
rect 1751 -3081 2071 -3039
<< properties >>
string FIXED_BBOX -2049 -3080 1511 3080
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 17 l 30 val 1.037k carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
