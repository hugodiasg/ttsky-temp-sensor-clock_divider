magic
tech sky130A
magscale 1 2
timestamp 1729294469
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 3 21 643 203
rect 28 -17 62 21
<< scnmos >>
rect 82 47 112 177
rect 168 47 198 177
rect 254 47 284 177
rect 362 47 392 177
rect 448 47 478 177
rect 534 47 564 177
<< scpmoshvt >>
rect 82 297 112 497
rect 168 297 198 497
rect 254 297 284 497
rect 354 297 384 497
rect 448 297 478 497
rect 534 297 564 497
<< ndiff >>
rect 29 165 82 177
rect 29 131 37 165
rect 71 131 82 165
rect 29 97 82 131
rect 29 63 37 97
rect 71 63 82 97
rect 29 47 82 63
rect 112 93 168 177
rect 112 59 123 93
rect 157 59 168 93
rect 112 47 168 59
rect 198 165 254 177
rect 198 131 209 165
rect 243 131 254 165
rect 198 97 254 131
rect 198 63 209 97
rect 243 63 254 97
rect 198 47 254 63
rect 284 93 362 177
rect 284 59 305 93
rect 339 59 362 93
rect 284 47 362 59
rect 392 165 448 177
rect 392 131 403 165
rect 437 131 448 165
rect 392 97 448 131
rect 392 63 403 97
rect 437 63 448 97
rect 392 47 448 63
rect 478 169 534 177
rect 478 135 489 169
rect 523 135 534 169
rect 478 47 534 135
rect 564 103 617 177
rect 564 69 575 103
rect 609 69 617 103
rect 564 47 617 69
<< pdiff >>
rect 29 485 82 497
rect 29 451 37 485
rect 71 451 82 485
rect 29 407 82 451
rect 29 373 37 407
rect 71 373 82 407
rect 29 297 82 373
rect 112 477 168 497
rect 112 443 123 477
rect 157 443 168 477
rect 112 407 168 443
rect 112 373 123 407
rect 157 373 168 407
rect 112 297 168 373
rect 198 409 254 497
rect 198 375 209 409
rect 243 375 254 409
rect 198 297 254 375
rect 284 477 354 497
rect 284 443 305 477
rect 339 443 354 477
rect 284 297 354 443
rect 384 485 448 497
rect 384 451 398 485
rect 432 451 448 485
rect 384 297 448 451
rect 478 435 534 497
rect 478 401 489 435
rect 523 401 534 435
rect 478 343 534 401
rect 478 309 489 343
rect 523 309 534 343
rect 478 297 534 309
rect 564 446 617 497
rect 564 412 575 446
rect 609 412 617 446
rect 564 364 617 412
rect 564 330 575 364
rect 609 330 617 364
rect 564 297 617 330
<< ndiffc >>
rect 37 131 71 165
rect 37 63 71 97
rect 123 59 157 93
rect 209 131 243 165
rect 209 63 243 97
rect 305 59 339 93
rect 403 131 437 165
rect 403 63 437 97
rect 489 135 523 169
rect 575 69 609 103
<< pdiffc >>
rect 37 451 71 485
rect 37 373 71 407
rect 123 443 157 477
rect 123 373 157 407
rect 209 375 243 409
rect 305 443 339 477
rect 398 451 432 485
rect 489 401 523 435
rect 489 309 523 343
rect 575 412 609 446
rect 575 330 609 364
<< poly >>
rect 82 497 112 523
rect 168 497 198 523
rect 254 497 284 523
rect 354 497 384 523
rect 448 497 478 523
rect 534 497 564 523
rect 82 261 112 297
rect 168 265 198 297
rect 254 265 284 297
rect 354 265 384 297
rect 24 249 112 261
rect 24 215 40 249
rect 74 215 112 249
rect 24 192 112 215
rect 154 249 284 265
rect 154 215 164 249
rect 198 215 233 249
rect 267 215 284 249
rect 154 199 284 215
rect 340 249 406 265
rect 340 215 356 249
rect 390 215 406 249
rect 340 199 406 215
rect 448 233 478 297
rect 534 265 564 297
rect 534 249 622 265
rect 534 233 576 249
rect 448 215 576 233
rect 610 215 622 249
rect 448 199 622 215
rect 82 177 112 192
rect 168 177 198 199
rect 254 177 284 199
rect 362 177 392 199
rect 448 192 564 199
rect 448 177 478 192
rect 534 177 564 192
rect 82 21 112 47
rect 168 21 198 47
rect 254 21 284 47
rect 362 21 392 47
rect 448 21 478 47
rect 534 21 564 47
<< polycont >>
rect 40 215 74 249
rect 164 215 198 249
rect 233 215 267 249
rect 356 215 390 249
rect 576 215 610 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 21 485 87 527
rect 21 451 37 485
rect 71 451 87 485
rect 21 407 87 451
rect 21 373 37 407
rect 71 373 87 407
rect 21 357 87 373
rect 121 477 343 493
rect 121 443 123 477
rect 157 459 305 477
rect 157 443 165 459
rect 121 407 165 443
rect 339 443 343 477
rect 305 427 343 443
rect 382 485 448 527
rect 382 451 398 485
rect 432 451 448 485
rect 382 435 448 451
rect 482 435 529 493
rect 121 373 123 407
rect 157 373 165 407
rect 121 357 165 373
rect 199 409 259 425
rect 199 375 209 409
rect 243 393 259 409
rect 482 401 489 435
rect 523 401 529 435
rect 482 393 529 401
rect 243 375 529 393
rect 199 357 529 375
rect 487 343 529 357
rect 24 289 419 323
rect 24 249 90 289
rect 24 215 40 249
rect 74 215 90 249
rect 124 249 284 255
rect 124 215 164 249
rect 198 215 233 249
rect 267 215 284 249
rect 320 249 419 289
rect 320 215 356 249
rect 390 215 419 249
rect 487 309 489 343
rect 523 309 529 343
rect 563 446 625 527
rect 563 412 575 446
rect 609 412 625 446
rect 563 364 625 412
rect 563 330 575 364
rect 609 330 625 364
rect 563 314 625 330
rect 24 211 90 215
rect 21 165 453 177
rect 21 131 37 165
rect 71 143 209 165
rect 71 131 87 143
rect 21 97 87 131
rect 193 131 209 143
rect 243 143 403 165
rect 243 131 259 143
rect 21 63 37 97
rect 71 63 87 97
rect 21 51 87 63
rect 123 93 157 109
rect 123 17 157 59
rect 193 97 259 131
rect 387 131 403 143
rect 437 131 453 165
rect 193 63 209 97
rect 243 63 259 97
rect 193 51 259 63
rect 305 93 339 109
rect 305 17 339 59
rect 387 97 453 131
rect 487 169 529 309
rect 487 135 489 169
rect 523 135 529 169
rect 563 249 626 280
rect 563 215 576 249
rect 610 215 626 249
rect 563 153 626 215
rect 487 119 529 135
rect 387 63 403 97
rect 437 85 453 97
rect 563 103 625 119
rect 563 85 575 103
rect 437 69 575 85
rect 609 69 625 103
rect 437 63 625 69
rect 387 51 625 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel locali s 580 153 614 187 0 FreeSans 200 0 0 0 B1
port 4 nsew
flabel locali s 488 357 522 391 0 FreeSans 200 0 0 0 Y
port 6 nsew
flabel locali s 396 357 430 391 0 FreeSans 200 0 0 0 Y
port 6 nsew
flabel locali s 304 357 338 391 0 FreeSans 200 0 0 0 Y
port 6 nsew
flabel locali s 212 221 246 255 0 FreeSans 200 0 0 0 A2
port 7 nsew
flabel locali s 212 357 246 391 0 FreeSans 200 0 0 0 Y
port 6 nsew
flabel locali s 28 289 62 323 0 FreeSans 200 0 0 0 A1
port 5 nsew
flabel locali s 28 221 62 255 0 FreeSans 200 0 0 0 A1
port 5 nsew
flabel locali s 580 221 614 255 0 FreeSans 200 0 0 0 B1
port 4 nsew
flabel metal1 s 28 -17 62 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 28 527 62 561 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 28 527 62 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew
flabel pwell s 28 -17 62 17 0 FreeSans 200 0 0 0 VNB
port 9 nsew
rlabel comment s 0 0 0 0 4 o21ai_2
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_END 257156
string GDS_FILE clock_divider.gds
string GDS_START 250712
string path 0.000 0.000 3.220 0.000 
<< end >>
