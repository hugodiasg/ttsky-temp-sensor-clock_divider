magic
tech sky130A
magscale 1 2
timestamp 1700762700
<< nwell >>
rect -581 -1600 581 1600
<< pmos >>
rect -487 -1500 -287 1500
rect -229 -1500 -29 1500
rect 29 -1500 229 1500
rect 287 -1500 487 1500
<< pdiff >>
rect -545 1488 -487 1500
rect -545 -1488 -533 1488
rect -499 -1488 -487 1488
rect -545 -1500 -487 -1488
rect -287 1488 -229 1500
rect -287 -1488 -275 1488
rect -241 -1488 -229 1488
rect -287 -1500 -229 -1488
rect -29 1488 29 1500
rect -29 -1488 -17 1488
rect 17 -1488 29 1488
rect -29 -1500 29 -1488
rect 229 1488 287 1500
rect 229 -1488 241 1488
rect 275 -1488 287 1488
rect 229 -1500 287 -1488
rect 487 1488 545 1500
rect 487 -1488 499 1488
rect 533 -1488 545 1488
rect 487 -1500 545 -1488
<< pdiffc >>
rect -533 -1488 -499 1488
rect -275 -1488 -241 1488
rect -17 -1488 17 1488
rect 241 -1488 275 1488
rect 499 -1488 533 1488
<< poly >>
rect -487 1581 -287 1597
rect -487 1547 -471 1581
rect -303 1547 -287 1581
rect -487 1500 -287 1547
rect -229 1581 -29 1597
rect -229 1547 -213 1581
rect -45 1547 -29 1581
rect -229 1500 -29 1547
rect 29 1581 229 1597
rect 29 1547 45 1581
rect 213 1547 229 1581
rect 29 1500 229 1547
rect 287 1581 487 1597
rect 287 1547 303 1581
rect 471 1547 487 1581
rect 287 1500 487 1547
rect -487 -1547 -287 -1500
rect -487 -1581 -471 -1547
rect -303 -1581 -287 -1547
rect -487 -1597 -287 -1581
rect -229 -1547 -29 -1500
rect -229 -1581 -213 -1547
rect -45 -1581 -29 -1547
rect -229 -1597 -29 -1581
rect 29 -1547 229 -1500
rect 29 -1581 45 -1547
rect 213 -1581 229 -1547
rect 29 -1597 229 -1581
rect 287 -1547 487 -1500
rect 287 -1581 303 -1547
rect 471 -1581 487 -1547
rect 287 -1597 487 -1581
<< polycont >>
rect -471 1547 -303 1581
rect -213 1547 -45 1581
rect 45 1547 213 1581
rect 303 1547 471 1581
rect -471 -1581 -303 -1547
rect -213 -1581 -45 -1547
rect 45 -1581 213 -1547
rect 303 -1581 471 -1547
<< locali >>
rect -487 1547 -471 1581
rect -303 1547 -287 1581
rect -229 1547 -213 1581
rect -45 1547 -29 1581
rect 29 1547 45 1581
rect 213 1547 229 1581
rect 287 1547 303 1581
rect 471 1547 487 1581
rect -533 1488 -499 1504
rect -533 -1504 -499 -1488
rect -275 1488 -241 1504
rect -275 -1504 -241 -1488
rect -17 1488 17 1504
rect -17 -1504 17 -1488
rect 241 1488 275 1504
rect 241 -1504 275 -1488
rect 499 1488 533 1504
rect 499 -1504 533 -1488
rect -487 -1581 -471 -1547
rect -303 -1581 -287 -1547
rect -229 -1581 -213 -1547
rect -45 -1581 -29 -1547
rect 29 -1581 45 -1547
rect 213 -1581 229 -1547
rect 287 -1581 303 -1547
rect 471 -1581 487 -1547
<< viali >>
rect -533 -17 -499 1471
rect -275 -1471 -241 17
rect -17 -17 17 1471
rect 241 -1471 275 17
rect 499 -17 533 1471
<< metal1 >>
rect -539 1471 -493 1483
rect -539 -17 -533 1471
rect -499 -17 -493 1471
rect -23 1471 23 1483
rect -539 -29 -493 -17
rect -281 17 -235 29
rect -281 -1471 -275 17
rect -241 -1471 -235 17
rect -23 -17 -17 1471
rect 17 -17 23 1471
rect 493 1471 539 1483
rect -23 -29 23 -17
rect 235 17 281 29
rect -281 -1483 -235 -1471
rect 235 -1471 241 17
rect 275 -1471 281 17
rect 493 -17 499 1471
rect 533 -17 539 1471
rect 493 -29 539 -17
rect 235 -1483 281 -1471
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 15.0 l 1.0 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc +50 viadrn -50 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
