magic
tech sky130A
timestamp 1701394307
<< pwell >>
rect -1598 -1605 1598 1605
<< nmos >>
rect -1500 -1500 1500 1500
<< ndiff >>
rect -1529 1494 -1500 1500
rect -1529 -1494 -1523 1494
rect -1506 -1494 -1500 1494
rect -1529 -1500 -1500 -1494
rect 1500 1494 1529 1500
rect 1500 -1494 1506 1494
rect 1523 -1494 1529 1494
rect 1500 -1500 1529 -1494
<< ndiffc >>
rect -1523 -1494 -1506 1494
rect 1506 -1494 1523 1494
<< psubdiff >>
rect -1580 1570 -1532 1587
rect 1532 1570 1580 1587
rect -1580 1539 -1563 1570
rect 1563 1539 1580 1570
rect -1580 -1570 -1563 -1539
rect 1563 -1570 1580 -1539
rect -1580 -1587 -1532 -1570
rect 1532 -1587 1580 -1570
<< psubdiffcont >>
rect -1532 1570 1532 1587
rect -1580 -1539 -1563 1539
rect 1563 -1539 1580 1539
rect -1532 -1587 1532 -1570
<< poly >>
rect -1500 1536 1500 1544
rect -1500 1519 -1492 1536
rect 1492 1519 1500 1536
rect -1500 1500 1500 1519
rect -1500 -1519 1500 -1500
rect -1500 -1536 -1492 -1519
rect 1492 -1536 1500 -1519
rect -1500 -1544 1500 -1536
<< polycont >>
rect -1492 1519 1492 1536
rect -1492 -1536 1492 -1519
<< locali >>
rect -1580 1570 -1532 1587
rect 1532 1570 1580 1587
rect -1580 1539 -1563 1570
rect 1563 1539 1580 1570
rect -1500 1519 -1492 1536
rect 1492 1519 1500 1536
rect -1523 1494 -1506 1502
rect -1523 -1502 -1506 -1494
rect 1506 1494 1523 1502
rect 1506 -1502 1523 -1494
rect -1500 -1536 -1492 -1519
rect 1492 -1536 1500 -1519
rect -1580 -1570 -1563 -1539
rect 1563 -1570 1580 -1539
rect -1580 -1587 -1532 -1570
rect 1532 -1587 1580 -1570
<< viali >>
rect -1492 1519 1492 1536
rect -1523 -1494 -1506 1494
rect 1506 -1494 1523 1494
rect -1492 -1536 1492 -1519
<< metal1 >>
rect -1498 1536 1498 1539
rect -1498 1519 -1492 1536
rect 1492 1519 1498 1536
rect -1498 1516 1498 1519
rect -1526 1494 -1503 1500
rect -1526 -1494 -1523 1494
rect -1506 -1494 -1503 1494
rect -1526 -1500 -1503 -1494
rect 1503 1494 1526 1500
rect 1503 -1494 1506 1494
rect 1523 -1494 1526 1494
rect 1503 -1500 1526 -1494
rect -1498 -1519 1498 -1516
rect -1498 -1536 -1492 -1519
rect 1492 -1536 1498 -1519
rect -1498 -1539 1498 -1536
<< properties >>
string FIXED_BBOX -1571 -1578 1571 1578
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 30 l 30 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
