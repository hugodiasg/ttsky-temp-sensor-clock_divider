magic
tech sky130A
timestamp 1701394307
<< pwell >>
rect -848 -1105 848 1105
<< nmos >>
rect -750 -1000 750 1000
<< ndiff >>
rect -779 994 -750 1000
rect -779 -994 -773 994
rect -756 -994 -750 994
rect -779 -1000 -750 -994
rect 750 994 779 1000
rect 750 -994 756 994
rect 773 -994 779 994
rect 750 -1000 779 -994
<< ndiffc >>
rect -773 -994 -756 994
rect 756 -994 773 994
<< psubdiff >>
rect -830 1070 -782 1087
rect 782 1070 830 1087
rect -830 1039 -813 1070
rect 813 1039 830 1070
rect -830 -1070 -813 -1039
rect 813 -1070 830 -1039
rect -830 -1087 -782 -1070
rect 782 -1087 830 -1070
<< psubdiffcont >>
rect -782 1070 782 1087
rect -830 -1039 -813 1039
rect 813 -1039 830 1039
rect -782 -1087 782 -1070
<< poly >>
rect -750 1036 750 1044
rect -750 1019 -742 1036
rect 742 1019 750 1036
rect -750 1000 750 1019
rect -750 -1019 750 -1000
rect -750 -1036 -742 -1019
rect 742 -1036 750 -1019
rect -750 -1044 750 -1036
<< polycont >>
rect -742 1019 742 1036
rect -742 -1036 742 -1019
<< locali >>
rect -830 1070 -782 1087
rect 782 1070 830 1087
rect -830 1039 -813 1070
rect 813 1039 830 1070
rect -750 1019 -742 1036
rect 742 1019 750 1036
rect -773 994 -756 1002
rect -773 -1002 -756 -994
rect 756 994 773 1002
rect 756 -1002 773 -994
rect -750 -1036 -742 -1019
rect 742 -1036 750 -1019
rect -830 -1070 -813 -1039
rect 813 -1070 830 -1039
rect -830 -1087 -782 -1070
rect 782 -1087 830 -1070
<< viali >>
rect -742 1019 742 1036
rect -773 -994 -756 994
rect 756 -994 773 994
rect -742 -1036 742 -1019
<< metal1 >>
rect -748 1036 748 1039
rect -748 1019 -742 1036
rect 742 1019 748 1036
rect -748 1016 748 1019
rect -776 994 -753 1000
rect -776 -994 -773 994
rect -756 -994 -753 994
rect -776 -1000 -753 -994
rect 753 994 776 1000
rect 753 -994 756 994
rect 773 -994 776 994
rect 753 -1000 776 -994
rect -748 -1019 748 -1016
rect -748 -1036 -742 -1019
rect 742 -1036 748 -1019
rect -748 -1039 748 -1036
<< properties >>
string FIXED_BBOX -821 -1078 821 1078
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 20 l 15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
