magic
tech sky130A
magscale 1 2
timestamp 1700703435
<< error_p >>
rect -229 328 -169 334
rect 169 328 229 334
rect -294 274 -275 308
rect -229 286 -164 328
rect 164 286 229 328
rect -229 274 -17 286
rect 17 274 229 286
rect -260 252 -164 274
rect -54 252 54 274
rect 164 252 260 274
rect -260 240 260 252
rect -260 212 -241 240
rect -275 178 -241 212
rect -260 -220 -241 178
rect -226 178 -172 240
rect -30 188 -29 189
rect -17 188 17 210
rect 29 188 30 189
rect -29 187 -28 188
rect -17 182 37 188
rect 84 182 122 210
rect 226 190 260 240
rect -226 -178 -214 178
rect -94 172 122 182
rect 214 178 260 190
rect -94 138 -84 172
rect -29 138 29 172
rect 84 138 122 172
rect -94 128 -17 138
rect 17 128 94 138
rect -18 100 -17 101
rect 17 100 37 128
rect -17 99 -16 100
rect 16 99 17 100
rect -157 88 -101 99
rect 101 88 157 99
rect -146 -77 -135 88
rect -112 -77 -101 88
rect -146 -88 -101 -77
rect 112 -77 123 88
rect 146 -77 157 88
rect 112 -88 157 -77
rect -17 -100 -16 -99
rect 16 -100 17 -99
rect -18 -101 -17 -100
rect 17 -128 37 -100
rect 84 -128 122 -100
rect -94 -138 -17 -128
rect 17 -138 122 -128
rect -94 -172 -84 -138
rect -29 -172 29 -138
rect 84 -172 122 -138
rect -226 -186 -172 -178
rect -94 -182 94 -172
rect 226 -178 238 178
rect 252 -178 260 178
rect -226 -220 -164 -186
rect -28 -187 37 -182
rect 226 -186 260 -178
rect -29 -188 37 -187
rect -30 -189 -29 -188
rect 29 -189 30 -188
rect -260 -228 -164 -220
rect 164 -228 260 -186
rect -260 -240 -17 -228
rect 17 -240 260 -228
rect -260 -262 -164 -240
rect -54 -262 54 -240
rect 164 -262 260 -240
rect -260 -274 260 -262
rect 275 -274 294 308
rect -229 -334 -169 -274
rect 169 -334 229 -274
<< pwell >>
rect -425 -710 425 710
<< nmos >>
rect -229 274 -29 500
rect 29 274 229 500
rect -226 188 -29 240
rect 29 188 226 240
rect -226 172 -17 188
rect 17 172 226 188
rect -226 138 -84 172
rect 84 138 226 172
rect -226 100 -17 138
rect 17 100 226 138
rect -226 88 226 100
rect -226 -88 -146 88
rect -112 -88 112 88
rect 146 -88 226 88
rect -226 -100 226 -88
rect -226 -138 -17 -100
rect 17 -138 226 -100
rect -226 -172 -84 -138
rect 84 -172 226 -138
rect -226 -188 -17 -172
rect 17 -188 226 -172
rect -226 -240 -29 -188
rect 29 -240 226 -188
rect -229 -500 -29 -274
rect 29 -500 229 -274
<< ndiff >>
rect -287 488 -229 500
rect -287 -488 -275 488
rect -241 274 -229 488
rect -29 488 29 500
rect -29 274 -17 488
rect 17 274 29 488
rect 229 488 287 500
rect 229 274 241 488
rect -29 188 -17 240
rect 17 188 29 240
rect -29 -240 -17 -188
rect 17 -240 29 -188
rect -241 -488 -229 -274
rect -287 -500 -229 -488
rect -29 -488 -17 -274
rect 17 -488 29 -274
rect -29 -500 29 -488
rect 229 -488 241 -274
rect 275 -488 287 488
rect 229 -500 287 -488
<< ndiffc >>
rect -275 274 -241 488
rect -17 274 17 488
rect 241 274 275 488
rect -275 -274 -260 274
rect -17 188 17 240
rect -146 -88 -112 88
rect 112 -88 146 88
rect -17 -240 17 -188
rect 260 -274 275 274
rect -275 -488 -241 -274
rect -17 -488 17 -274
rect 241 -488 275 -274
<< psubdiff >>
rect -389 640 -293 674
rect 293 640 389 674
rect -389 578 -355 640
rect 355 578 389 640
rect -260 240 -164 274
rect 164 240 260 274
rect -260 178 -226 240
rect 226 178 260 240
rect -260 -240 -226 -178
rect 226 -240 260 -178
rect -260 -274 -164 -240
rect 164 -274 260 -240
rect -389 -640 -355 -578
rect 355 -640 389 -578
rect -389 -674 -293 -640
rect 293 -674 389 -640
<< psubdiffcont >>
rect -293 640 293 674
rect -389 -578 -355 578
rect -164 240 164 274
rect -260 -178 -226 178
rect 226 -178 260 178
rect -164 -274 164 -240
rect 355 -578 389 578
rect -293 -674 293 -640
<< poly >>
rect -229 572 -29 588
rect -229 538 -213 572
rect -45 538 -29 572
rect -229 500 -29 538
rect 29 572 229 588
rect 29 538 45 572
rect 213 538 229 572
rect 29 500 229 538
rect -17 172 17 188
rect -17 100 17 138
rect -17 -138 17 -100
rect -17 -188 17 -172
rect -229 -538 -29 -500
rect -229 -572 -213 -538
rect -45 -572 -29 -538
rect -229 -588 -29 -572
rect 29 -538 229 -500
rect 29 -572 45 -538
rect 213 -572 229 -538
rect 29 -588 229 -572
<< polycont >>
rect -213 538 -45 572
rect 45 538 213 572
rect -84 138 84 172
rect -84 -172 84 -138
rect -213 -572 -45 -538
rect 45 -572 213 -538
<< locali >>
rect -389 640 -293 674
rect 293 640 389 674
rect -389 578 -355 640
rect 355 578 389 640
rect -229 538 -213 572
rect -45 538 -29 572
rect 29 538 45 572
rect 213 538 229 572
rect -275 488 -241 504
rect -17 488 17 504
rect 241 488 275 504
rect -241 240 -164 274
rect 164 240 241 274
rect -241 178 -226 240
rect 226 178 241 240
rect -100 138 -84 172
rect 84 138 100 172
rect -146 88 -112 104
rect -146 -104 -112 -88
rect 112 88 146 104
rect 112 -104 146 -88
rect -100 -172 -84 -138
rect 84 -172 100 -138
rect -241 -240 -226 -178
rect 226 -240 241 -178
rect -241 -274 -164 -240
rect 164 -274 241 -240
rect -275 -504 -241 -488
rect -17 -504 17 -488
rect 241 -504 275 -488
rect -229 -572 -213 -538
rect -45 -572 -29 -538
rect 29 -572 45 -538
rect 213 -572 229 -538
rect -389 -640 -355 -578
rect 355 -640 389 -578
rect -389 -674 -293 -640
rect 293 -674 389 -640
<< viali >>
rect -213 538 -45 572
rect 45 538 213 572
rect -275 274 -241 488
rect -17 274 17 488
rect 241 274 275 488
rect -275 -274 -260 274
rect -260 178 -241 274
rect -17 240 17 274
rect -260 -178 -241 178
rect -17 188 17 240
rect -17 172 17 188
rect 241 178 260 274
rect -84 138 84 172
rect -146 -88 -112 88
rect -17 -138 17 138
rect 112 -88 146 88
rect -84 -172 84 -138
rect -260 -274 -241 -178
rect -17 -188 17 -172
rect -17 -240 17 -188
rect 241 -178 260 178
rect -17 -274 17 -240
rect 241 -274 260 -178
rect 260 -274 275 274
rect -275 -488 -241 -274
rect -17 -488 17 -274
rect 241 -488 275 -274
rect -213 -572 -45 -538
rect 45 -572 213 -538
<< metal1 >>
rect -225 572 -33 578
rect -225 538 -213 572
rect -45 538 -33 572
rect -225 532 -33 538
rect 33 572 225 578
rect 33 538 45 572
rect 213 538 225 572
rect 33 532 225 538
rect -281 488 -235 500
rect -281 -488 -275 488
rect -241 -488 -235 488
rect -23 488 23 500
rect -23 178 -17 488
rect -96 172 -17 178
rect 17 178 23 488
rect 235 488 281 500
rect 17 172 96 178
rect -96 138 -84 172
rect 84 138 96 172
rect -96 132 -17 138
rect -152 88 -106 100
rect -152 -88 -146 88
rect -112 -88 -106 88
rect -152 -100 -106 -88
rect -23 -132 -17 132
rect -96 -138 -17 -132
rect 17 132 96 138
rect 17 -132 23 132
rect 106 88 152 100
rect 106 -88 112 88
rect 146 -88 152 88
rect 106 -100 152 -88
rect 17 -138 96 -132
rect -96 -172 -84 -138
rect 84 -172 96 -138
rect -96 -178 -17 -172
rect -281 -500 -235 -488
rect -23 -488 -17 -178
rect 17 -178 96 -172
rect 17 -488 23 -178
rect -23 -500 23 -488
rect 235 -488 241 488
rect 275 -488 281 488
rect 235 -500 281 -488
rect -225 -538 -33 -532
rect -225 -572 -213 -538
rect -45 -572 -33 -538
rect -225 -578 -33 -572
rect 33 -538 225 -532
rect 33 -572 45 -538
rect 213 -572 225 -538
rect 33 -578 225 -572
<< properties >>
string FIXED_BBOX -243 -257 243 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
