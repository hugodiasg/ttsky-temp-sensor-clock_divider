magic
tech sky130A
magscale 1 2
timestamp 1700708449
<< metal4 >>
rect -3349 839 3349 880
rect -3349 -839 3093 839
rect 3329 -839 3349 839
rect -3349 -880 3349 -839
<< via4 >>
rect 3093 -839 3329 839
<< mimcap2 >>
rect -3269 760 2731 800
rect -3269 -760 -3229 760
rect 2691 -760 2731 760
rect -3269 -800 2731 -760
<< mimcap2contact >>
rect -3229 -760 2691 760
<< metal5 >>
rect 3051 839 3371 881
rect -3253 760 2715 784
rect -3253 -760 -3229 760
rect 2691 -760 2715 760
rect -3253 -784 2715 -760
rect 3051 -839 3093 839
rect 3329 -839 3371 839
rect 3051 -881 3371 -839
<< properties >>
string FIXED_BBOX -3349 -880 2811 880
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 30 l 8 val 494.44 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
