magic
tech sky130A
magscale 1 2
timestamp 1699929776
<< nmos >>
rect -100 527 100 727
rect -100 109 100 309
rect -100 -309 100 -109
rect -100 -727 100 -527
<< ndiff >>
rect -158 715 -100 727
rect -158 539 -146 715
rect -112 539 -100 715
rect -158 527 -100 539
rect 100 715 158 727
rect 100 539 112 715
rect 146 539 158 715
rect 100 527 158 539
rect -158 297 -100 309
rect -158 121 -146 297
rect -112 121 -100 297
rect -158 109 -100 121
rect 100 297 158 309
rect 100 121 112 297
rect 146 121 158 297
rect 100 109 158 121
rect -158 -121 -100 -109
rect -158 -297 -146 -121
rect -112 -297 -100 -121
rect -158 -309 -100 -297
rect 100 -121 158 -109
rect 100 -297 112 -121
rect 146 -297 158 -121
rect 100 -309 158 -297
rect -158 -539 -100 -527
rect -158 -715 -146 -539
rect -112 -715 -100 -539
rect -158 -727 -100 -715
rect 100 -539 158 -527
rect 100 -715 112 -539
rect 146 -715 158 -539
rect 100 -727 158 -715
<< ndiffc >>
rect -146 539 -112 715
rect 112 539 146 715
rect -146 121 -112 297
rect 112 121 146 297
rect -146 -297 -112 -121
rect 112 -297 146 -121
rect -146 -715 -112 -539
rect 112 -715 146 -539
<< poly >>
rect -100 799 100 815
rect -100 765 -84 799
rect 84 765 100 799
rect -100 727 100 765
rect -100 489 100 527
rect -100 455 -84 489
rect 84 455 100 489
rect -100 439 100 455
rect -100 381 100 397
rect -100 347 -84 381
rect 84 347 100 381
rect -100 309 100 347
rect -100 71 100 109
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -109 100 -71
rect -100 -347 100 -309
rect -100 -381 -84 -347
rect 84 -381 100 -347
rect -100 -397 100 -381
rect -100 -455 100 -439
rect -100 -489 -84 -455
rect 84 -489 100 -455
rect -100 -527 100 -489
rect -100 -765 100 -727
rect -100 -799 -84 -765
rect 84 -799 100 -765
rect -100 -815 100 -799
<< polycont >>
rect -84 765 84 799
rect -84 455 84 489
rect -84 347 84 381
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -381 84 -347
rect -84 -489 84 -455
rect -84 -799 84 -765
<< locali >>
rect -100 765 -84 799
rect 84 765 100 799
rect -146 715 -112 731
rect -146 523 -112 539
rect 112 715 146 731
rect 112 523 146 539
rect -100 455 -84 489
rect 84 455 100 489
rect -100 347 -84 381
rect 84 347 100 381
rect -146 297 -112 313
rect -146 105 -112 121
rect 112 297 146 313
rect 112 105 146 121
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -121 -112 -105
rect -146 -313 -112 -297
rect 112 -121 146 -105
rect 112 -313 146 -297
rect -100 -381 -84 -347
rect 84 -381 100 -347
rect -100 -489 -84 -455
rect 84 -489 100 -455
rect -146 -539 -112 -523
rect -146 -731 -112 -715
rect 112 -539 146 -523
rect 112 -731 146 -715
rect -100 -799 -84 -765
rect 84 -799 100 -765
<< viali >>
rect -84 765 84 799
rect -146 539 -112 715
rect 112 539 146 715
rect -84 455 84 489
rect -84 347 84 381
rect -146 121 -112 297
rect 112 121 146 297
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -297 -112 -121
rect 112 -297 146 -121
rect -84 -381 84 -347
rect -84 -489 84 -455
rect -146 -715 -112 -539
rect 112 -715 146 -539
rect -84 -799 84 -765
<< metal1 >>
rect -96 799 96 805
rect -96 765 -84 799
rect 84 765 96 799
rect -96 759 96 765
rect -152 715 -106 727
rect -152 539 -146 715
rect -112 539 -106 715
rect -152 527 -106 539
rect 106 715 152 727
rect 106 539 112 715
rect 146 539 152 715
rect 106 527 152 539
rect -96 489 96 495
rect -96 455 -84 489
rect 84 455 96 489
rect -96 449 96 455
rect -96 381 96 387
rect -96 347 -84 381
rect 84 347 96 381
rect -96 341 96 347
rect -152 297 -106 309
rect -152 121 -146 297
rect -112 121 -106 297
rect -152 109 -106 121
rect 106 297 152 309
rect 106 121 112 297
rect 146 121 152 297
rect 106 109 152 121
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -121 -106 -109
rect -152 -297 -146 -121
rect -112 -297 -106 -121
rect -152 -309 -106 -297
rect 106 -121 152 -109
rect 106 -297 112 -121
rect 146 -297 152 -121
rect 106 -309 152 -297
rect -96 -347 96 -341
rect -96 -381 -84 -347
rect 84 -381 96 -347
rect -96 -387 96 -381
rect -96 -455 96 -449
rect -96 -489 -84 -455
rect 84 -489 96 -455
rect -96 -495 96 -489
rect -152 -539 -106 -527
rect -152 -715 -146 -539
rect -112 -715 -106 -539
rect -152 -727 -106 -715
rect 106 -539 152 -527
rect 106 -715 112 -539
rect 146 -715 152 -539
rect 106 -727 152 -715
rect -96 -765 96 -759
rect -96 -799 -84 -765
rect 84 -799 96 -765
rect -96 -805 96 -799
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 1.0 m 4 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
