magic
tech sky130A
magscale 1 2
timestamp 1700703435
<< metal4 >>
rect -2549 2439 2549 2480
rect -2549 -2439 2293 2439
rect 2529 -2439 2549 2439
rect -2549 -2480 2549 -2439
<< via4 >>
rect 2293 -2439 2529 2439
<< mimcap2 >>
rect -2469 2360 1931 2400
rect -2469 -2360 -2429 2360
rect 1891 -2360 1931 2360
rect -2469 -2400 1931 -2360
<< mimcap2contact >>
rect -2429 -2360 1891 2360
<< metal5 >>
rect 2251 2439 2571 2481
rect -2453 2360 1915 2384
rect -2453 -2360 -2429 2360
rect 1891 -2360 1915 2360
rect -2453 -2384 1915 -2360
rect 2251 -2439 2293 2439
rect 2529 -2439 2571 2439
rect 2251 -2481 2571 -2439
<< properties >>
string FIXED_BBOX -2549 -2480 2011 2480
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 22 l 24 val 1.073k carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
