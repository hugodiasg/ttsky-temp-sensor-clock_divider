magic
tech sky130A
timestamp 1699933188
<< pwell >>
rect -1098 -555 1098 555
<< nmos >>
rect -1000 -450 1000 450
<< ndiff >>
rect -1029 444 -1000 450
rect -1029 -444 -1023 444
rect -1006 -444 -1000 444
rect -1029 -450 -1000 -444
rect 1000 444 1029 450
rect 1000 -444 1006 444
rect 1023 -444 1029 444
rect 1000 -450 1029 -444
<< ndiffc >>
rect -1023 -444 -1006 444
rect 1006 -444 1023 444
<< psubdiff >>
rect -1080 520 -1032 537
rect 1032 520 1080 537
rect -1080 489 -1063 520
rect 1063 489 1080 520
rect -1080 -520 -1063 -489
rect 1063 -520 1080 -489
rect -1080 -537 -1032 -520
rect 1032 -537 1080 -520
<< psubdiffcont >>
rect -1032 520 1032 537
rect -1080 -489 -1063 489
rect 1063 -489 1080 489
rect -1032 -537 1032 -520
<< poly >>
rect -1000 486 1000 494
rect -1000 469 -992 486
rect 992 469 1000 486
rect -1000 450 1000 469
rect -1000 -469 1000 -450
rect -1000 -486 -992 -469
rect 992 -486 1000 -469
rect -1000 -494 1000 -486
<< polycont >>
rect -992 469 992 486
rect -992 -486 992 -469
<< locali >>
rect -1080 520 -1032 537
rect 1032 520 1080 537
rect -1080 489 -1063 520
rect 1063 489 1080 520
rect -1000 469 -992 486
rect 992 469 1000 486
rect -1023 444 -1006 452
rect -1023 -452 -1006 -444
rect 1006 444 1023 452
rect 1006 -452 1023 -444
rect -1000 -486 -992 -469
rect 992 -486 1000 -469
rect -1080 -520 -1063 -489
rect 1063 -520 1080 -489
rect -1080 -537 -1032 -520
rect 1032 -537 1080 -520
<< viali >>
rect -992 469 992 486
rect -1023 -444 -1006 444
rect 1006 -444 1023 444
rect -992 -486 992 -469
<< metal1 >>
rect -998 486 998 489
rect -998 469 -992 486
rect 992 469 998 486
rect -998 466 998 469
rect -1026 444 -1003 450
rect -1026 -444 -1023 444
rect -1006 -444 -1003 444
rect -1026 -450 -1003 -444
rect 1003 444 1026 450
rect 1003 -444 1006 444
rect 1023 -444 1026 444
rect 1003 -450 1026 -444
rect -998 -469 998 -466
rect -998 -486 -992 -469
rect 992 -486 998 -469
rect -998 -489 998 -486
<< properties >>
string FIXED_BBOX -1071 -528 1071 528
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 9 l 20 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
