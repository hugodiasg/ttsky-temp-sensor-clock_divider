magic
tech sky130A
magscale 1 2
timestamp 1699935153
<< nwell >>
rect -453 1127 3573 2793
rect -493 -193 2733 873
<< pwell >>
rect -660 -2340 2732 -420
<< psubdiff >>
rect -624 -490 -528 -456
rect 2600 -490 2696 -456
rect -624 -552 -590 -490
rect -624 -2270 -590 -2208
rect 2662 -552 2696 -490
rect 2662 -2270 2696 -2208
rect -624 -2304 -528 -2270
rect 2600 -2304 2696 -2270
<< nsubdiff >>
rect -417 2723 -357 2757
rect 3477 2723 3537 2757
rect -417 2697 -383 2723
rect -417 1197 -383 1223
rect 3503 2697 3537 2723
rect 3503 1197 3537 1223
rect -417 1163 -357 1197
rect 3477 1163 3537 1197
rect -457 803 -397 837
rect 2637 803 2697 837
rect -457 777 -423 803
rect -457 -123 -423 -97
rect 2663 777 2697 803
rect 2663 -123 2697 -97
rect -457 -157 -397 -123
rect 2637 -157 2697 -123
<< psubdiffcont >>
rect -528 -490 2600 -456
rect -624 -2208 -590 -552
rect 2662 -2208 2696 -552
rect -528 -2304 2600 -2270
<< nsubdiffcont >>
rect -357 2723 3477 2757
rect -417 1223 -383 2697
rect 3503 1223 3537 2697
rect -357 1163 3477 1197
rect -397 803 2637 837
rect -457 -97 -423 777
rect 2663 -97 2697 777
rect -397 -157 2637 -123
<< locali >>
rect -417 2723 -357 2757
rect 3477 2723 3537 2757
rect -417 2697 -383 2723
rect -417 1197 -383 1223
rect 3503 2697 3537 2723
rect 3503 1197 3537 1223
rect -417 1163 -357 1197
rect 3477 1163 3537 1197
rect -457 803 -397 837
rect 2637 803 2697 837
rect -457 777 -423 803
rect 2663 777 2697 803
rect -457 -123 -423 -97
rect 2663 -123 2697 -97
rect -457 -157 -397 -123
rect 2637 -157 2697 -123
rect -624 -490 -528 -456
rect 2600 -490 2696 -456
rect -624 -552 -590 -490
rect -624 -2270 -590 -2208
rect 2662 -552 2696 -490
rect 2662 -2270 2696 -2208
rect -624 -2304 -528 -2270
rect 2600 -2304 2696 -2270
<< viali >>
rect 180 2757 340 2760
rect 1300 2757 1460 2760
rect 2080 2757 2240 2760
rect 3000 2757 3160 2760
rect 180 2723 340 2757
rect 1300 2723 1460 2757
rect 2080 2723 2240 2757
rect 3000 2723 3160 2757
rect 180 2720 340 2723
rect 1300 2720 1460 2723
rect 2080 2720 2240 2723
rect 3000 2720 3160 2723
rect 2620 440 2663 540
rect 2663 440 2697 540
rect 2697 440 2700 540
rect -440 -2270 -220 -2260
rect 440 -2270 660 -2260
rect 1360 -2270 1580 -2260
rect 2200 -2270 2420 -2260
rect -440 -2300 -220 -2270
rect 440 -2300 660 -2270
rect 1360 -2300 1580 -2270
rect 2200 -2300 2420 -2270
<< metal1 >>
rect -340 2900 3580 3000
rect -350 2800 -340 2900
rect -260 2800 940 2900
rect 1060 2800 3380 2900
rect 3480 2800 3580 2900
rect 180 2766 340 2800
rect 1300 2766 1460 2800
rect 2080 2766 2240 2800
rect 3000 2766 3160 2800
rect 168 2760 352 2766
rect 168 2720 180 2760
rect 340 2720 352 2760
rect 168 2714 352 2720
rect 1288 2760 1472 2766
rect 1288 2720 1300 2760
rect 1460 2720 1472 2760
rect 1288 2714 1472 2720
rect 2068 2760 2252 2766
rect 2068 2720 2080 2760
rect 2240 2720 2252 2760
rect 2068 2714 2252 2720
rect 2988 2760 3172 2766
rect 2988 2720 3000 2760
rect 3160 2720 3172 2760
rect 2988 2714 3172 2720
rect 1160 2560 1380 2580
rect 1140 2460 1380 2560
rect 3100 2540 3320 2560
rect 3060 2460 3320 2540
rect 930 2340 940 2460
rect 1060 2340 1540 2460
rect 2920 2340 3380 2460
rect 3480 2340 3490 2460
rect 2920 2320 3360 2340
rect 1690 2080 1700 2300
rect 1780 2080 1790 2300
rect 1860 2240 2720 2260
rect 1860 2120 2620 2240
rect 2720 2120 2730 2240
rect 1540 2000 1960 2040
rect 1950 1980 1960 2000
rect 2060 1980 2070 2040
rect -220 1800 -20 1880
rect -350 1720 -340 1800
rect -260 1720 400 1800
rect 1000 1700 1700 1800
rect 1780 1700 1840 1800
rect 2160 1680 2260 1780
rect 2360 1680 2720 1780
rect 100 1360 660 1520
rect 740 1400 3380 1500
rect 100 1340 180 1360
rect 160 1300 180 1340
rect 280 1300 1760 1360
rect 1950 1300 1960 1360
rect 2060 1320 2920 1360
rect 3120 1320 3300 1400
rect 2060 1300 2070 1320
rect 3380 1040 3580 1060
rect 1950 920 1960 1040
rect 2060 920 3580 1040
rect 1960 900 3580 920
rect 3380 860 3580 900
rect -280 540 -20 660
rect 2300 540 2520 660
rect 2614 540 2706 552
rect 3380 540 3580 600
rect -300 440 2620 540
rect 2740 440 3580 540
rect 2614 428 2706 440
rect 3380 400 3580 440
rect 80 280 2180 300
rect 80 80 1960 280
rect 2040 80 2180 280
rect 80 60 2180 80
rect 1370 -80 1380 -20
rect 1440 -80 2260 -20
rect 2360 -80 2370 -20
rect -130 -260 -120 -180
rect -60 -200 520 -180
rect -60 -260 180 -200
rect 280 -260 520 -200
rect 580 -260 590 -180
rect 630 -220 640 -140
rect 700 -220 1280 -140
rect 1340 -220 1960 -140
rect 2060 -220 2070 -140
rect 2030 -420 2040 -340
rect 2100 -420 2260 -340
rect 2340 -420 2350 -340
rect -500 -2260 -180 -530
rect 2010 -540 2020 -520
rect -60 -580 2020 -540
rect 2100 -580 2110 -520
rect 2360 -560 2480 -550
rect 2200 -600 2480 -560
rect -130 -810 -120 -630
rect -60 -810 -50 -630
rect 150 -830 160 -630
rect 300 -830 310 -630
rect 510 -810 520 -630
rect 580 -810 590 -630
rect 630 -810 640 -650
rect 700 -810 710 -650
rect 920 -670 1060 -630
rect 910 -810 920 -670
rect 1020 -810 1060 -670
rect 920 -830 1060 -810
rect 1250 -820 1260 -640
rect 1320 -820 1330 -640
rect 1370 -830 1380 -630
rect 1460 -830 1470 -630
rect 1680 -650 1820 -630
rect 1670 -810 1680 -650
rect 1800 -810 1820 -650
rect 2010 -830 2020 -650
rect 2080 -830 2090 -650
rect 0 -1000 100 -860
rect 360 -1020 460 -880
rect 740 -1020 840 -880
rect 1140 -1020 1240 -880
rect 1520 -1020 1620 -880
rect 1880 -1020 1980 -880
rect -130 -1250 -120 -1050
rect -60 -1250 -50 -1050
rect 150 -1250 160 -1050
rect 300 -1250 310 -1050
rect 510 -1230 520 -1050
rect 580 -1230 590 -1050
rect 630 -1230 640 -1070
rect 700 -1230 710 -1070
rect 920 -1090 1060 -1050
rect 920 -1230 940 -1090
rect 1040 -1230 1060 -1090
rect 920 -1250 1060 -1230
rect 1250 -1240 1260 -1060
rect 1320 -1240 1330 -1060
rect 1390 -1250 1400 -1050
rect 1480 -1250 1490 -1050
rect 1680 -1070 1820 -1050
rect 1670 -1230 1680 -1070
rect 1800 -1230 1820 -1070
rect 2030 -1230 2040 -1050
rect 2100 -1230 2110 -1050
rect 0 -1420 100 -1280
rect 360 -1420 460 -1278
rect 740 -1420 840 -1278
rect 1140 -1420 1240 -1278
rect 1520 -1420 1620 -1278
rect 1880 -1420 1980 -1278
rect -130 -1650 -120 -1470
rect -60 -1650 -50 -1470
rect 150 -1670 160 -1470
rect 300 -1670 310 -1470
rect 510 -1650 520 -1470
rect 580 -1650 590 -1470
rect 630 -1650 640 -1490
rect 700 -1650 710 -1490
rect 920 -1510 1060 -1470
rect 920 -1650 940 -1510
rect 1040 -1650 1060 -1510
rect 920 -1670 1060 -1650
rect 1250 -1660 1260 -1480
rect 1320 -1660 1330 -1480
rect 1390 -1650 1400 -1470
rect 1460 -1650 1470 -1470
rect 1680 -1490 1820 -1470
rect 1670 -1650 1680 -1490
rect 1800 -1650 1820 -1490
rect 2030 -1650 2040 -1470
rect 2100 -1650 2110 -1470
rect 0 -1840 100 -1700
rect 360 -1840 460 -1696
rect 740 -1840 840 -1696
rect 1140 -1840 1240 -1696
rect 1520 -1840 1620 -1696
rect 1880 -1840 1980 -1696
rect -130 -2070 -120 -1890
rect -60 -2070 -50 -1890
rect 150 -2070 160 -1890
rect 300 -2070 310 -1890
rect 510 -2070 520 -1890
rect 580 -2070 590 -1890
rect 630 -2070 640 -1910
rect 700 -2070 710 -1910
rect 920 -1930 1060 -1890
rect 920 -2070 940 -1930
rect 1040 -2070 1060 -1930
rect 920 -2090 1060 -2070
rect 1250 -2080 1260 -1900
rect 1320 -2080 1330 -1900
rect 1390 -2070 1400 -1890
rect 1460 -2070 1470 -1890
rect 1680 -1910 1820 -1890
rect 1670 -2070 1680 -1910
rect 1800 -2070 1820 -1910
rect 2030 -2070 2040 -1890
rect 2100 -2070 2110 -1890
rect -500 -2300 -440 -2260
rect -220 -2290 -180 -2260
rect 428 -2260 672 -2254
rect 428 -2290 440 -2260
rect -220 -2300 440 -2290
rect 660 -2290 672 -2260
rect 1348 -2260 1592 -2254
rect 1348 -2290 1360 -2260
rect 660 -2300 920 -2290
rect -500 -2310 920 -2300
rect -500 -2410 180 -2310
rect 280 -2410 920 -2310
rect -500 -2430 920 -2410
rect 1040 -2300 1360 -2290
rect 1580 -2290 1592 -2260
rect 2160 -2260 2480 -600
rect 2160 -2290 2200 -2260
rect 1580 -2300 1680 -2290
rect 1040 -2430 1680 -2300
rect 1820 -2300 2200 -2290
rect 2420 -2300 2480 -2260
rect 1820 -2430 2480 -2300
rect -500 -2500 2480 -2430
<< via1 >>
rect -340 2800 -260 2900
rect 940 2800 1060 2900
rect 3380 2800 3480 2900
rect 940 2340 1060 2460
rect 3380 2340 3480 2460
rect 1700 2080 1780 2300
rect 2620 2120 2720 2240
rect 1960 1980 2060 2040
rect -340 1720 -260 1800
rect 1700 1700 1780 1800
rect 2260 1680 2360 1780
rect 180 1300 280 1360
rect 1960 1300 2060 1360
rect 1960 920 2060 1040
rect 2620 440 2700 540
rect 2700 440 2740 540
rect 1960 80 2040 280
rect 1380 -80 1440 -20
rect 2260 -80 2360 -20
rect -120 -260 -60 -180
rect 180 -260 280 -200
rect 520 -260 580 -180
rect 640 -220 700 -140
rect 1280 -220 1340 -140
rect 1960 -220 2060 -140
rect 2040 -420 2100 -340
rect 2260 -420 2340 -340
rect 2020 -580 2100 -520
rect -120 -810 -60 -630
rect 160 -830 300 -630
rect 520 -810 580 -630
rect 640 -810 700 -650
rect 920 -810 1020 -670
rect 1260 -820 1320 -640
rect 1380 -830 1460 -630
rect 1680 -810 1800 -650
rect 2020 -830 2080 -650
rect -120 -1250 -60 -1050
rect 160 -1250 300 -1050
rect 520 -1230 580 -1050
rect 640 -1230 700 -1070
rect 940 -1230 1040 -1090
rect 1260 -1240 1320 -1060
rect 1400 -1250 1480 -1050
rect 1680 -1230 1800 -1070
rect 2040 -1230 2100 -1050
rect -120 -1650 -60 -1470
rect 160 -1670 300 -1470
rect 520 -1650 580 -1470
rect 640 -1650 700 -1490
rect 940 -1650 1040 -1510
rect 1260 -1660 1320 -1480
rect 1400 -1650 1460 -1470
rect 1680 -1650 1800 -1490
rect 2040 -1650 2100 -1470
rect -120 -2070 -60 -1890
rect 160 -2070 300 -1890
rect 520 -2070 580 -1890
rect 640 -2070 700 -1910
rect 940 -2070 1040 -1930
rect 1260 -2080 1320 -1900
rect 1400 -2070 1460 -1890
rect 1680 -2070 1800 -1910
rect 2040 -2070 2100 -1890
rect 180 -2410 280 -2310
rect 920 -2430 1040 -2290
rect 1680 -2430 1820 -2290
<< metal2 >>
rect -340 2900 -260 2910
rect -340 1800 -260 2800
rect 940 2900 1060 2910
rect 940 2460 1060 2800
rect 940 2330 1060 2340
rect 3380 2900 3480 2910
rect 3380 2460 3480 2800
rect 3380 2330 3480 2340
rect -340 1710 -260 1720
rect 1700 2300 1780 2310
rect 1700 1800 1780 2080
rect 2620 2240 2740 2260
rect 2720 2120 2740 2240
rect 1700 1690 1780 1700
rect 1960 2040 2060 2050
rect 180 1360 280 1370
rect -120 -180 -60 -170
rect -120 -630 -60 -260
rect 180 -200 280 1300
rect 1960 1360 2060 1980
rect 1960 1040 2060 1300
rect 1960 280 2060 920
rect 2040 80 2060 280
rect 1380 -20 1440 -10
rect 640 -140 700 -130
rect 180 -270 280 -260
rect 520 -180 580 -170
rect -120 -1050 -60 -810
rect -120 -1470 -60 -1250
rect -120 -1890 -60 -1650
rect -120 -2090 -60 -2070
rect 160 -630 300 -620
rect 160 -1050 300 -830
rect 160 -1470 300 -1250
rect 160 -1890 300 -1670
rect 160 -2310 300 -2070
rect 520 -630 580 -260
rect 520 -1050 580 -810
rect 520 -1470 580 -1230
rect 520 -1890 580 -1650
rect 520 -2090 580 -2070
rect 640 -650 700 -220
rect 1280 -140 1340 -130
rect 1280 -630 1340 -220
rect 1260 -640 1340 -630
rect 640 -1070 700 -810
rect 640 -1490 700 -1230
rect 640 -1910 700 -1650
rect 640 -2090 700 -2070
rect 920 -670 1040 -650
rect 1020 -810 1040 -670
rect 920 -1090 1040 -810
rect 1320 -820 1340 -640
rect 1260 -830 1340 -820
rect 1280 -1050 1340 -830
rect 920 -1230 940 -1090
rect 920 -1510 1040 -1230
rect 1260 -1060 1340 -1050
rect 1320 -1240 1340 -1060
rect 1260 -1250 1340 -1240
rect 1280 -1470 1340 -1250
rect 920 -1650 940 -1510
rect 920 -1930 1040 -1650
rect 1260 -1480 1340 -1470
rect 1320 -1660 1340 -1480
rect 1260 -1670 1340 -1660
rect 1280 -1890 1340 -1670
rect 920 -2070 940 -1930
rect 160 -2410 180 -2310
rect 280 -2410 300 -2310
rect 160 -2430 300 -2410
rect 920 -2290 1040 -2070
rect 1260 -1900 1340 -1890
rect 1320 -2080 1340 -1900
rect 1260 -2090 1340 -2080
rect 1380 -620 1440 -80
rect 1960 -140 2060 80
rect 1960 -230 2060 -220
rect 2260 1780 2360 1790
rect 2260 -20 2360 1680
rect 2620 540 2740 2120
rect 2620 430 2740 440
rect 2260 -110 2360 -80
rect 2040 -340 2100 -330
rect 2040 -510 2100 -420
rect 2260 -340 2340 -110
rect 2260 -430 2340 -420
rect 2020 -520 2100 -510
rect 2020 -590 2100 -580
rect 1380 -630 1460 -620
rect 1380 -840 1460 -830
rect 1680 -650 1820 -630
rect 2040 -640 2100 -590
rect 1800 -810 1820 -650
rect 1380 -1040 1440 -840
rect 1380 -1050 1480 -1040
rect 1380 -1250 1400 -1050
rect 1380 -1260 1480 -1250
rect 1680 -1070 1820 -810
rect 2020 -650 2100 -640
rect 2080 -830 2100 -650
rect 2020 -840 2100 -830
rect 1800 -1230 1820 -1070
rect 1380 -1460 1440 -1260
rect 1380 -1470 1460 -1460
rect 1380 -1650 1400 -1470
rect 1380 -1660 1460 -1650
rect 1680 -1490 1820 -1230
rect 1800 -1650 1820 -1490
rect 1380 -1880 1440 -1660
rect 1380 -1890 1460 -1880
rect 1380 -2070 1400 -1890
rect 1380 -2080 1460 -2070
rect 1680 -1910 1820 -1650
rect 1800 -2070 1820 -1910
rect 1380 -2150 1440 -2080
rect 920 -2440 1040 -2430
rect 1680 -2290 1820 -2070
rect 2040 -1050 2100 -840
rect 2040 -1470 2100 -1230
rect 2040 -1890 2100 -1650
rect 2040 -2130 2100 -2070
rect 1680 -2440 1820 -2430
use sky130_fd_pr__nfet_01v8_9VJR3B  sky130_fd_pr__nfet_01v8_9VJR3B_0
timestamp 1699929776
transform 1 0 -342 0 1 -1355
box -158 -815 158 815
use sky130_fd_pr__nfet_01v8_9VJR3B  sky130_fd_pr__nfet_01v8_9VJR3B_1
timestamp 1699929776
transform 1 0 38 0 1 -1355
box -158 -815 158 815
use sky130_fd_pr__nfet_01v8_9VJR3B  sky130_fd_pr__nfet_01v8_9VJR3B_2
timestamp 1699929776
transform 1 0 418 0 1 -1355
box -158 -815 158 815
use sky130_fd_pr__nfet_01v8_9VJR3B  sky130_fd_pr__nfet_01v8_9VJR3B_3
timestamp 1699929776
transform 1 0 798 0 1 -1355
box -158 -815 158 815
use sky130_fd_pr__nfet_01v8_9VJR3B  sky130_fd_pr__nfet_01v8_9VJR3B_4
timestamp 1699929776
transform 1 0 1178 0 1 -1355
box -158 -815 158 815
use sky130_fd_pr__nfet_01v8_9VJR3B  sky130_fd_pr__nfet_01v8_9VJR3B_5
timestamp 1699929776
transform 1 0 1558 0 1 -1355
box -158 -815 158 815
use sky130_fd_pr__nfet_01v8_9VJR3B  sky130_fd_pr__nfet_01v8_9VJR3B_6
timestamp 1699929776
transform 1 0 2318 0 1 -1355
box -158 -815 158 815
use sky130_fd_pr__nfet_01v8_9VJR3B  sky130_fd_pr__nfet_01v8_9VJR3B_7
timestamp 1699929776
transform 1 0 1938 0 1 -1355
box -158 -815 158 815
use sky130_fd_pr__pfet_01v8_FRXWNM  sky130_fd_pr__pfet_01v8_FRXWNM_0
timestamp 1699932112
transform 1 0 -126 0 1 1600
box -194 -300 194 300
use sky130_fd_pr__pfet_01v8_FRXWNM  sky130_fd_pr__pfet_01v8_FRXWNM_1
timestamp 1699932112
transform 1 0 1254 0 1 2280
box -194 -300 194 300
use sky130_fd_pr__pfet_01v8_FRXWNM  sky130_fd_pr__pfet_01v8_FRXWNM_2
timestamp 1699932112
transform 1 0 3194 0 1 2280
box -194 -300 194 300
use sky130_fd_pr__pfet_01v8_FRXWNM  sky130_fd_pr__pfet_01v8_FRXWNM_3
timestamp 1699932112
transform 1 0 -146 0 1 360
box -194 -300 194 300
use sky130_fd_pr__pfet_01v8_FRXWNM  sky130_fd_pr__pfet_01v8_FRXWNM_4
timestamp 1699932112
transform 1 0 2414 0 1 360
box -194 -300 194 300
use sky130_fd_pr__pfet_01v8_FVXEPM  sky130_fd_pr__pfet_01v8_FVXEPM_0
timestamp 1699932112
transform 1 0 3214 0 1 1600
box -194 -300 194 300
use sky130_fd_pr__pfet_01v8_YAEUFM  sky130_fd_pr__pfet_01v8_YAEUFM_0
timestamp 1699932112
transform 1 0 1137 0 1 360
box -1097 -300 1097 300
use sky130_fd_pr__pfet_01v8_YAWWFM  sky130_fd_pr__pfet_01v8_YAWWFM_0
timestamp 1699932112
transform 1 0 1281 0 1 1600
box -581 -300 581 300
use sky130_fd_pr__pfet_01v8_YAWWFM  sky130_fd_pr__pfet_01v8_YAWWFM_1
timestamp 1699932112
transform 1 0 2441 0 1 1600
box -581 -300 581 300
use sky130_fd_pr__pfet_01v8_FVTXNM  XP1
timestamp 1699932112
transform 1 0 383 0 1 1600
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_3HGYVM  XP3
timestamp 1699929776
transform 1 0 1634 0 1 2280
box -194 -300 194 300
use sky130_fd_pr__pfet_01v8_SKTYVM  XP4
timestamp 1699929776
transform 1 0 2414 0 1 2280
box -594 -300 594 300
<< labels >>
flabel metal1 -180 2800 20 3000 0 FreeSans 256 0 0 0 vd
port 0 nsew
flabel metal1 -500 -2500 -300 -2300 0 FreeSans 256 0 0 0 gnd
port 3 nsew
flabel metal1 3380 400 3580 600 0 FreeSans 256 0 0 0 vts
port 1 nsew
flabel metal1 3380 860 3580 1060 0 FreeSans 256 0 0 0 vtd
port 2 nsew
flabel metal2 200 1080 220 1100 0 FreeSans 800 0 0 0 a
flabel metal2 1720 1940 1740 1960 0 FreeSans 800 0 0 0 d
flabel metal1 1840 1440 1860 1480 0 FreeSans 800 0 0 0 c
flabel metal2 2300 -280 2300 -260 0 FreeSans 800 0 0 0 b
<< end >>
