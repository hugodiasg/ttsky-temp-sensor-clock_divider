magic
tech sky130A
magscale 1 2
timestamp 1723762448
<< error_p >>
rect -29 381 29 387
rect -29 347 -17 381
rect -29 341 29 347
rect -29 -347 29 -341
rect -29 -381 -17 -347
rect -29 -387 29 -381
<< nwell >>
rect -211 -519 211 519
<< pmos >>
rect -15 -300 15 300
<< pdiff >>
rect -73 288 -15 300
rect -73 -288 -61 288
rect -27 -288 -15 288
rect -73 -300 -15 -288
rect 15 288 73 300
rect 15 -288 27 288
rect 61 -288 73 288
rect 15 -300 73 -288
<< pdiffc >>
rect -61 -288 -27 288
rect 27 -288 61 288
<< nsubdiff >>
rect -175 449 -79 483
rect 79 449 175 483
rect -175 387 -141 449
rect 141 387 175 449
rect -175 -449 -141 -387
rect 141 -449 175 -387
rect -175 -483 -79 -449
rect 79 -483 175 -449
<< nsubdiffcont >>
rect -79 449 79 483
rect -175 -387 -141 387
rect 141 -387 175 387
rect -79 -483 79 -449
<< poly >>
rect -33 381 33 397
rect -33 347 -17 381
rect 17 347 33 381
rect -33 331 33 347
rect -15 300 15 331
rect -15 -331 15 -300
rect -33 -347 33 -331
rect -33 -381 -17 -347
rect 17 -381 33 -347
rect -33 -397 33 -381
<< polycont >>
rect -17 347 17 381
rect -17 -381 17 -347
<< locali >>
rect -175 449 -79 483
rect 79 449 175 483
rect -175 387 -141 449
rect 141 387 175 449
rect -33 347 -17 381
rect 17 347 33 381
rect -61 288 -27 304
rect -61 -304 -27 -288
rect 27 288 61 304
rect 27 -304 61 -288
rect -33 -381 -17 -347
rect 17 -381 33 -347
rect -175 -449 -141 -387
rect 141 -449 175 -387
rect -175 -483 -79 -449
rect 79 -483 175 -449
<< viali >>
rect -17 347 17 381
rect -61 -288 -27 288
rect 27 -288 61 288
rect -17 -381 17 -347
<< metal1 >>
rect -29 381 29 387
rect -29 347 -17 381
rect 17 347 29 381
rect -29 341 29 347
rect -67 288 -21 300
rect -67 -288 -61 288
rect -27 -288 -21 288
rect -67 -300 -21 -288
rect 21 288 67 300
rect 21 -288 27 288
rect 61 -288 67 288
rect 21 -300 67 -288
rect -29 -347 29 -341
rect -29 -381 -17 -347
rect 17 -381 29 -347
rect -29 -387 29 -381
<< properties >>
string FIXED_BBOX -158 -466 158 466
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 3.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
