magic
tech sky130A
magscale 1 2
timestamp 1700703435
<< pwell >>
rect -1225 -310 1225 310
<< nmos >>
rect -1029 -100 -29 100
rect 29 -100 1029 100
<< ndiff >>
rect -1087 88 -1029 100
rect -1087 -88 -1075 88
rect -1041 -88 -1029 88
rect -1087 -100 -1029 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 1029 88 1087 100
rect 1029 -88 1041 88
rect 1075 -88 1087 88
rect 1029 -100 1087 -88
<< ndiffc >>
rect -1075 -88 -1041 88
rect -17 -88 17 88
rect 1041 -88 1075 88
<< psubdiff >>
rect -1189 240 -1093 274
rect 1093 240 1189 274
rect -1189 178 -1155 240
rect 1155 178 1189 240
rect -1189 -240 -1155 -178
rect 1155 -240 1189 -178
rect -1189 -274 -1093 -240
rect 1093 -274 1189 -240
<< psubdiffcont >>
rect -1093 240 1093 274
rect -1189 -178 -1155 178
rect 1155 -178 1189 178
rect -1093 -274 1093 -240
<< poly >>
rect -1029 172 -29 188
rect -1029 138 -1013 172
rect -45 138 -29 172
rect -1029 100 -29 138
rect 29 172 1029 188
rect 29 138 45 172
rect 1013 138 1029 172
rect 29 100 1029 138
rect -1029 -138 -29 -100
rect -1029 -172 -1013 -138
rect -45 -172 -29 -138
rect -1029 -188 -29 -172
rect 29 -138 1029 -100
rect 29 -172 45 -138
rect 1013 -172 1029 -138
rect 29 -188 1029 -172
<< polycont >>
rect -1013 138 -45 172
rect 45 138 1013 172
rect -1013 -172 -45 -138
rect 45 -172 1013 -138
<< locali >>
rect -1189 240 -1093 274
rect 1093 240 1189 274
rect -1189 178 -1155 240
rect 1155 178 1189 240
rect -1029 138 -1013 172
rect -45 138 -29 172
rect 29 138 45 172
rect 1013 138 1029 172
rect -1075 88 -1041 104
rect -1075 -104 -1041 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 1041 88 1075 104
rect 1041 -104 1075 -88
rect -1029 -172 -1013 -138
rect -45 -172 -29 -138
rect 29 -172 45 -138
rect 1013 -172 1029 -138
rect -1189 -240 -1155 -178
rect 1155 -240 1189 -178
rect -1189 -274 -1093 -240
rect 1093 -274 1189 -240
<< viali >>
rect -1013 138 -45 172
rect 45 138 1013 172
rect -1075 -88 -1041 88
rect -17 -88 17 88
rect 1041 -88 1075 88
rect -1013 -172 -45 -138
rect 45 -172 1013 -138
<< metal1 >>
rect -1025 172 -33 178
rect -1025 138 -1013 172
rect -45 138 -33 172
rect -1025 132 -33 138
rect 33 172 1025 178
rect 33 138 45 172
rect 1013 138 1025 172
rect 33 132 1025 138
rect -1081 88 -1035 100
rect -1081 -88 -1075 88
rect -1041 -88 -1035 88
rect -1081 -100 -1035 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 1035 88 1081 100
rect 1035 -88 1041 88
rect 1075 -88 1081 88
rect 1035 -100 1081 -88
rect -1025 -138 -33 -132
rect -1025 -172 -1013 -138
rect -45 -172 -33 -138
rect -1025 -178 -33 -172
rect 33 -138 1025 -132
rect 33 -172 45 -138
rect 1013 -172 1025 -138
rect 33 -178 1025 -172
<< properties >>
string FIXED_BBOX -1172 -257 1172 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 5 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
