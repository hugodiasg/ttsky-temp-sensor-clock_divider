magic
tech sky130A
magscale 1 2
timestamp 1707919911
<< metal3 >>
rect -3186 1512 3186 1540
rect -3186 -1512 3102 1512
rect 3166 -1512 3186 1512
rect -3186 -1540 3186 -1512
<< via3 >>
rect 3102 -1512 3166 1512
<< mimcap >>
rect -3146 1460 2854 1500
rect -3146 -1460 -3106 1460
rect 2814 -1460 2854 1460
rect -3146 -1500 2854 -1460
<< mimcapcontact >>
rect -3106 -1460 2814 1460
<< metal4 >>
rect 3086 1512 3182 1528
rect -3107 1460 2815 1461
rect -3107 -1460 -3106 1460
rect 2814 -1460 2815 1460
rect -3107 -1461 2815 -1460
rect 3086 -1512 3102 1512
rect 3166 -1512 3182 1512
rect 3086 -1528 3182 -1512
<< properties >>
string FIXED_BBOX -3186 -1540 2894 1540
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30 l 15 val 917.1 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
