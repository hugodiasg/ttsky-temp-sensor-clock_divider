magic
tech sky130A
magscale 1 2
timestamp 1700703435
<< metal4 >>
rect -2849 1539 2849 1580
rect -2849 -1539 2593 1539
rect 2829 -1539 2849 1539
rect -2849 -1580 2849 -1539
<< via4 >>
rect 2593 -1539 2829 1539
<< mimcap2 >>
rect -2769 1460 2231 1500
rect -2769 -1460 -2729 1460
rect 2191 -1460 2231 1460
rect -2769 -1500 2231 -1460
<< mimcap2contact >>
rect -2729 -1460 2191 1460
<< metal5 >>
rect 2551 1539 2871 1581
rect -2753 1460 2215 1484
rect -2753 -1460 -2729 1460
rect 2191 -1460 2215 1460
rect -2753 -1484 2215 -1460
rect 2551 -1539 2593 1539
rect 2829 -1539 2871 1539
rect 2551 -1581 2871 -1539
<< properties >>
string FIXED_BBOX -2849 -1580 2311 1580
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 25 l 15 val 765.2 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
