magic
tech sky130A
magscale 1 2
timestamp 1700747285
<< nmos >>
rect -1300 -900 1300 900
<< ndiff >>
rect -1358 888 -1300 900
rect -1358 -888 -1346 888
rect -1312 -888 -1300 888
rect -1358 -900 -1300 -888
rect 1300 888 1358 900
rect 1300 -888 1312 888
rect 1346 -888 1358 888
rect 1300 -900 1358 -888
<< ndiffc >>
rect -1346 -888 -1312 888
rect 1312 -888 1346 888
<< poly >>
rect -1300 972 1300 988
rect -1300 938 -1284 972
rect 1284 938 1300 972
rect -1300 900 1300 938
rect -1300 -938 1300 -900
rect -1300 -972 -1284 -938
rect 1284 -972 1300 -938
rect -1300 -988 1300 -972
<< polycont >>
rect -1284 938 1284 972
rect -1284 -972 1284 -938
<< locali >>
rect -1300 938 -1284 972
rect 1284 938 1300 972
rect -1346 888 -1312 904
rect -1346 -904 -1312 -888
rect 1312 888 1346 904
rect 1312 -904 1346 -888
rect -1300 -972 -1284 -938
rect 1284 -972 1300 -938
<< viali >>
rect -1284 938 1284 972
rect -1346 -871 -1312 17
rect 1312 -17 1346 871
rect -1284 -972 1284 -938
<< metal1 >>
rect -1296 972 1296 978
rect -1296 938 -1284 972
rect 1284 938 1296 972
rect -1296 932 1296 938
rect 1306 871 1352 883
rect -1352 17 -1306 29
rect -1352 -871 -1346 17
rect -1312 -871 -1306 17
rect 1306 -17 1312 871
rect 1346 -17 1352 871
rect 1306 -29 1352 -17
rect -1352 -883 -1306 -871
rect -1296 -938 1296 -932
rect -1296 -972 -1284 -938
rect 1284 -972 1296 -938
rect -1296 -978 1296 -972
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 9 l 13 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc -50 viadrn +50 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
