magic
tech sky130A
magscale 1 2
timestamp 1700703435
<< metal4 >>
rect -2549 2239 2549 2280
rect -2549 -2239 2293 2239
rect 2529 -2239 2549 2239
rect -2549 -2280 2549 -2239
<< via4 >>
rect 2293 -2239 2529 2239
<< mimcap2 >>
rect -2469 2160 1931 2200
rect -2469 -2160 -2429 2160
rect 1891 -2160 1931 2160
rect -2469 -2200 1931 -2160
<< mimcap2contact >>
rect -2429 -2160 1891 2160
<< metal5 >>
rect 2251 2239 2571 2281
rect -2453 2160 1915 2184
rect -2453 -2160 -2429 2160
rect 1891 -2160 1915 2160
rect -2453 -2184 1915 -2160
rect 2251 -2239 2293 2239
rect 2529 -2239 2571 2239
rect 2251 -2281 2571 -2239
<< properties >>
string FIXED_BBOX -2549 -2280 2011 2280
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 22 l 22 val 984.72 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
