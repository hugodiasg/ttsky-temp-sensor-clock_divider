magic
tech sky130A
magscale 1 2
timestamp 1738709249
<< metal1 >>
rect 10690 13140 10700 13480
rect 11000 13140 11010 13480
rect 10740 12900 10940 13140
rect 18940 12520 19140 12560
rect 18930 12260 18940 12520
rect 19160 12260 19170 12520
rect 2970 11780 2980 11940
rect 3160 11780 3170 11940
rect 18940 11680 19140 12260
rect 14030 10420 14040 10600
rect 14220 10420 14230 10600
rect 15060 10320 16100 10340
rect 15060 10140 15100 10320
rect 15280 10140 16100 10320
rect 6340 9520 7560 9540
rect 6340 9360 6660 9520
rect 6840 9360 7560 9520
rect 6340 9340 7560 9360
rect 7080 9160 7560 9180
rect 7080 8980 7100 9160
rect 7300 8980 7560 9160
rect 15700 7740 16100 7760
rect 15700 7600 15740 7740
rect 15860 7600 16100 7740
rect 15700 7560 16100 7600
rect 15380 7300 15400 7460
rect 15580 7300 15960 7460
rect 15380 7260 15960 7300
rect 14740 6940 14760 7120
rect 14920 6940 16100 7120
rect 14740 6920 16100 6940
rect 2430 6380 2440 6540
rect 2660 6380 2670 6540
rect 15390 6360 15400 6540
rect 15600 6360 16100 6560
rect 7350 5500 7360 5640
rect 7560 5500 7570 5640
<< via1 >>
rect 10700 13140 11000 13480
rect 18940 12260 19160 12520
rect 2980 11780 3160 11940
rect 14040 10420 14220 10600
rect 15100 10140 15280 10320
rect 6660 9360 6840 9520
rect 7100 8980 7300 9160
rect 15740 7600 15860 7740
rect 15400 7300 15580 7460
rect 14760 6940 14920 7120
rect 2440 6380 2660 6540
rect 15400 6360 15600 6540
rect 7360 5500 7560 5640
<< metal2 >>
rect 13360 41040 13520 41050
rect 7480 41020 7620 41030
rect 7480 40870 7620 40880
rect 10420 41020 10560 41030
rect 19240 41040 19400 41050
rect 13360 40930 13520 40940
rect 16280 41020 16440 41030
rect 10420 40850 10560 40860
rect 22200 41020 22320 41030
rect 28080 41020 28220 41030
rect 22200 40910 22320 40920
rect 25140 40980 25260 40990
rect 19240 40890 19400 40900
rect 28080 40910 28220 40920
rect 25140 40870 25260 40880
rect 16280 40830 16440 40840
rect 14740 16240 14940 16260
rect 14740 16060 14760 16240
rect 14920 16060 14940 16240
rect 10700 13480 11000 13490
rect 10700 13130 11000 13140
rect 2940 12300 3180 12310
rect 2940 12050 3180 12060
rect 2980 11940 3160 12050
rect 2980 11770 3160 11780
rect 14020 10600 14220 10620
rect 14020 10420 14040 10600
rect 6640 9520 6840 9540
rect 6640 9360 6660 9520
rect 2440 6540 2660 6550
rect 2440 6370 2660 6380
rect 2460 6190 2640 6370
rect 2440 6180 2680 6190
rect 2440 5910 2680 5920
rect 6640 2700 6840 9360
rect 7080 9170 7280 9180
rect 7080 9160 7300 9170
rect 7080 8980 7100 9160
rect 7080 8970 7300 8980
rect 7080 3180 7280 8970
rect 7360 5640 7560 5650
rect 7360 5350 7560 5500
rect 7360 5340 7580 5350
rect 7360 5090 7580 5100
rect 14020 3820 14220 10420
rect 14740 7120 14940 16060
rect 18940 14140 19160 14150
rect 15400 14080 15600 14100
rect 14740 6940 14760 7120
rect 14920 6940 14940 7120
rect 14740 6920 14940 6940
rect 15080 10320 15300 10340
rect 15080 10140 15100 10320
rect 15280 10140 15300 10320
rect 15080 4160 15300 10140
rect 15400 7460 15600 13900
rect 18940 12520 19160 13880
rect 18940 12250 19160 12260
rect 15740 7740 15860 7750
rect 15740 7590 15860 7600
rect 15580 7300 15600 7460
rect 15400 6540 15600 7300
rect 15400 6350 15600 6360
rect 16180 4890 16320 6180
rect 16160 4880 16340 4890
rect 16160 4630 16340 4640
rect 15260 3980 15300 4160
rect 15080 3950 15300 3980
rect 14020 3640 14040 3820
rect 14040 3630 14220 3640
rect 7080 2980 7280 3000
rect 6640 2540 6660 2700
rect 6640 2520 6840 2540
<< via2 >>
rect 7480 40880 7620 41020
rect 10420 40860 10560 41020
rect 13360 40940 13520 41040
rect 16280 40840 16440 41020
rect 19240 40900 19400 41040
rect 22200 40920 22320 41020
rect 25140 40880 25260 40980
rect 28080 40920 28220 41020
rect 14760 16060 14920 16240
rect 10700 13140 11000 13480
rect 2940 12060 3180 12300
rect 2440 5920 2680 6180
rect 7360 5100 7580 5340
rect 15400 13900 15600 14080
rect 18940 13880 19160 14140
rect 15740 7600 15860 7740
rect 16160 4640 16340 4880
rect 15080 3980 15260 4160
rect 14040 3640 14220 3820
rect 7080 3000 7280 3180
rect 6660 2540 6840 2700
<< metal3 >>
rect 4610 44640 4620 44780
rect 4740 44640 14940 44780
rect 15060 44640 15080 44780
rect 25150 44760 25270 44765
rect 25120 44660 25140 44760
rect 25260 44660 27080 44760
rect 25150 44635 25270 44660
rect 27070 44640 27080 44660
rect 27180 44640 27190 44760
rect 27610 44640 27620 44760
rect 27760 44640 28100 44760
rect 28200 44640 28210 44760
rect 22190 44400 22200 44520
rect 22320 44420 26540 44520
rect 26620 44420 26630 44520
rect 22320 44400 22330 44420
rect 22210 44395 22310 44400
rect 19250 44280 19390 44285
rect 19250 44120 19260 44280
rect 19400 44270 19410 44280
rect 19400 44260 26090 44270
rect 19400 44140 25980 44260
rect 26080 44140 26090 44260
rect 19400 44130 26090 44140
rect 19400 44120 19410 44130
rect 19250 44115 19390 44120
rect 16270 43820 16280 44000
rect 16440 43980 16450 44000
rect 16440 43820 25420 43980
rect 25540 43820 25560 43980
rect 16290 43815 16450 43820
rect 13370 43640 13530 43645
rect 13360 43500 13380 43640
rect 13500 43500 24840 43640
rect 24980 43500 25010 43640
rect 13370 43495 13530 43500
rect 10430 43340 10570 43345
rect 10400 43200 10440 43340
rect 10540 43200 24320 43340
rect 24440 43200 24450 43340
rect 10430 43195 10570 43200
rect 7470 43080 7650 43085
rect 7470 43060 23740 43080
rect 7470 42920 7480 43060
rect 7620 42920 23740 43060
rect 23900 42920 23910 43080
rect 7470 42915 7650 42920
rect 5830 42540 5840 42680
rect 6000 42660 6010 42680
rect 6000 42540 18800 42660
rect 18900 42540 18910 42660
rect 5850 42535 5990 42540
rect 5450 42140 5460 42280
rect 5620 42260 5630 42280
rect 5620 42140 28420 42260
rect 28540 42140 28550 42260
rect 5470 42135 5610 42140
rect 5050 41760 5060 41920
rect 5200 41919 5210 41920
rect 28710 41919 28720 41920
rect 5200 41760 28720 41919
rect 28860 41900 29720 41920
rect 28860 41760 29540 41900
rect 28720 41720 29540 41760
rect 29700 41720 29720 41900
rect 13350 41040 13530 41045
rect 7470 41020 7630 41025
rect 7470 40880 7480 41020
rect 7620 40880 7630 41020
rect 7470 40875 7630 40880
rect 10410 41020 10570 41025
rect 10410 40860 10420 41020
rect 10560 40860 10570 41020
rect 13350 40940 13360 41040
rect 13520 40940 13530 41040
rect 19230 41040 19410 41045
rect 13350 40935 13530 40940
rect 16270 41020 16450 41025
rect 10410 40855 10570 40860
rect 16270 40840 16280 41020
rect 16440 40840 16450 41020
rect 19230 40900 19240 41040
rect 19400 40900 19410 41040
rect 22190 41020 22330 41025
rect 22190 40920 22200 41020
rect 22320 40920 22330 41020
rect 28070 41020 28230 41025
rect 22190 40915 22330 40920
rect 25130 40980 25270 40985
rect 19230 40895 19410 40900
rect 25130 40880 25140 40980
rect 25260 40880 25270 40980
rect 28070 40920 28080 41020
rect 28220 40920 28230 41020
rect 28070 40915 28230 40920
rect 25130 40875 25270 40880
rect 16270 40835 16450 40840
rect 5850 36740 5990 36745
rect 5830 36600 5840 36740
rect 6000 36600 6010 36740
rect 5450 28720 5460 28860
rect 5620 28848 5630 28860
rect 5620 28728 5980 28848
rect 5620 28720 5630 28728
rect 5470 28715 5610 28720
rect 5050 20840 5060 20960
rect 5220 20840 6000 20960
rect 850 17440 860 17520
rect 820 17280 860 17440
rect 1140 17440 1150 17520
rect 1140 17420 25460 17440
rect 1140 17280 25280 17420
rect 25460 17280 25470 17420
rect 290 16960 300 17240
rect 520 17160 530 17240
rect 520 17000 26000 17160
rect 26120 17000 26140 17160
rect 520 16960 530 17000
rect 4590 16500 4600 16640
rect 4720 16630 4730 16640
rect 4720 16620 15870 16630
rect 4720 16500 15740 16620
rect 4610 16490 15740 16500
rect 15730 16480 15740 16490
rect 15860 16480 15870 16620
rect 14740 16240 29540 16260
rect 14740 16060 14760 16240
rect 14920 16080 29540 16240
rect 29700 16080 29720 16260
rect 14920 16060 29720 16080
rect 14750 16055 14930 16060
rect 18930 14140 19170 14145
rect 290 13860 300 14120
rect 520 14100 530 14120
rect 18930 14100 18940 14140
rect 520 14080 18940 14100
rect 520 13900 15400 14080
rect 15600 13900 18940 14080
rect 520 13880 18940 13900
rect 19160 13880 19170 14140
rect 520 13860 530 13880
rect 18930 13875 19170 13880
rect 270 13220 280 13560
rect 580 13480 590 13560
rect 10690 13480 11010 13485
rect 580 13280 10700 13480
rect 580 13220 590 13280
rect 10690 13140 10700 13280
rect 11000 13140 11010 13480
rect 10690 13135 11010 13140
rect 290 12080 300 12320
rect 600 12300 610 12320
rect 2930 12300 3190 12305
rect 600 12080 2940 12300
rect 2930 12060 2940 12080
rect 3180 12060 3190 12300
rect 2930 12055 3190 12060
rect 15730 7740 15870 7745
rect 15730 7600 15740 7740
rect 15860 7600 15870 7740
rect 15730 7595 15870 7600
rect 2430 6180 2690 6185
rect 870 5940 880 6180
rect 1160 6160 1170 6180
rect 2430 6160 2440 6180
rect 1160 5960 2440 6160
rect 1160 5940 1170 5960
rect 2430 5920 2440 5960
rect 2680 5920 2690 6180
rect 2430 5915 2690 5920
rect 860 5345 7560 5360
rect 860 5340 7590 5345
rect 860 5320 7360 5340
rect 860 5100 920 5320
rect 1140 5100 7360 5320
rect 7580 5100 7590 5340
rect 7350 5095 7590 5100
rect 830 4620 840 4900
rect 1140 4860 1150 4900
rect 16150 4880 16350 4885
rect 16150 4860 16160 4880
rect 1140 4640 16160 4860
rect 16340 4860 16350 4880
rect 16340 4640 16360 4860
rect 1140 4620 16360 4640
rect 15080 4165 30550 4170
rect 15070 4160 30550 4165
rect 15070 3980 15080 4160
rect 15260 4140 30550 4160
rect 15260 3980 30340 4140
rect 15070 3975 30340 3980
rect 15080 3960 30340 3975
rect 30520 3960 30550 4140
rect 15080 3950 30550 3960
rect 14020 3820 26500 3840
rect 14020 3640 14040 3820
rect 14220 3660 26500 3820
rect 26680 3660 26700 3840
rect 14220 3640 26700 3660
rect 14030 3635 14230 3640
rect 7070 3180 7290 3185
rect 7070 3000 7080 3180
rect 7280 3000 22620 3180
rect 22820 3000 22840 3180
rect 7070 2995 22840 3000
rect 7080 2980 22840 2995
rect 6640 2700 18940 2720
rect 6640 2540 6660 2700
rect 6840 2540 18760 2700
rect 18940 2540 18950 2700
rect 6640 2520 18940 2540
<< via3 >>
rect 4620 44640 4740 44780
rect 14940 44640 15060 44780
rect 25140 44660 25260 44760
rect 27080 44640 27180 44760
rect 27620 44640 27760 44760
rect 28100 44640 28200 44760
rect 22200 44400 22320 44520
rect 26540 44420 26620 44520
rect 19260 44120 19400 44280
rect 25980 44140 26080 44260
rect 16280 43820 16440 44000
rect 25420 43820 25540 43980
rect 13380 43500 13500 43640
rect 24840 43500 24980 43640
rect 10440 43200 10540 43340
rect 24320 43200 24440 43340
rect 7480 42920 7620 43060
rect 23740 42920 23900 43080
rect 5840 42540 6000 42680
rect 18800 42540 18900 42660
rect 5460 42140 5620 42280
rect 28420 42140 28540 42260
rect 5060 41760 5200 41920
rect 28720 41760 28860 41920
rect 29540 41720 29700 41900
rect 7480 40880 7620 41020
rect 10420 40860 10560 41020
rect 13360 40940 13520 41040
rect 16280 40840 16440 41020
rect 19240 40900 19400 41040
rect 22200 40920 22320 41020
rect 25140 40880 25260 40980
rect 28080 40920 28220 41020
rect 5840 36600 6000 36740
rect 5460 28720 5620 28860
rect 5060 20840 5220 20960
rect 860 17280 1140 17520
rect 25280 17280 25460 17420
rect 300 16960 520 17240
rect 26000 17000 26120 17160
rect 4600 16500 4720 16640
rect 15740 16480 15860 16620
rect 29540 16080 29700 16260
rect 300 13860 520 14120
rect 280 13220 580 13560
rect 300 12080 600 12320
rect 15740 7600 15860 7740
rect 880 5940 1160 6180
rect 920 5100 1140 5320
rect 840 4620 1140 4900
rect 30340 3960 30520 4140
rect 26500 3660 26680 3840
rect 22620 3000 22820 3180
rect 18760 2540 18940 2700
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44781 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 4619 44780 4741 44781
rect 14939 44780 15061 44781
rect 4610 44640 4620 44780
rect 4740 44640 4750 44780
rect 200 17240 600 44152
rect 200 16960 300 17240
rect 520 16960 600 17240
rect 200 14120 600 16960
rect 200 13860 300 14120
rect 520 13860 600 14120
rect 200 13560 600 13860
rect 200 13220 280 13560
rect 580 13220 600 13560
rect 200 12321 600 13220
rect 800 17520 1200 44152
rect 800 17280 860 17520
rect 1140 17280 1200 17520
rect 200 12320 601 12321
rect 200 12080 300 12320
rect 600 12080 601 12320
rect 200 12079 601 12080
rect 200 1000 600 12079
rect 800 6180 1200 17280
rect 4610 16641 4750 44640
rect 14939 44640 14940 44780
rect 15060 44640 15061 44780
rect 14939 44639 15061 44640
rect 16279 44000 16441 44001
rect 16279 43820 16280 44000
rect 16440 43820 16460 44000
rect 16279 43819 16460 43820
rect 13360 43640 13520 43660
rect 13360 43500 13380 43640
rect 13500 43500 13520 43640
rect 10420 43340 10560 43380
rect 10420 43200 10440 43340
rect 10540 43200 10560 43340
rect 7460 43060 7640 43120
rect 7460 42920 7480 43060
rect 7620 42920 7640 43060
rect 5839 42680 6001 42681
rect 5839 42540 5840 42680
rect 6000 42540 6001 42680
rect 5839 42539 6001 42540
rect 5460 42281 5620 42300
rect 5459 42280 5621 42281
rect 5459 42140 5460 42280
rect 5620 42140 5621 42280
rect 5459 42139 5621 42140
rect 5059 41920 5201 41921
rect 5059 41760 5060 41920
rect 5200 41919 5201 41920
rect 5200 41760 5220 41919
rect 5059 41759 5220 41760
rect 5061 20961 5220 41759
rect 5460 28861 5620 42139
rect 5840 36741 6000 42539
rect 7460 41020 7640 42920
rect 10420 41021 10560 43200
rect 13360 41041 13520 43500
rect 13359 41040 13521 41041
rect 7460 40880 7480 41020
rect 7620 40880 7640 41020
rect 7460 40860 7640 40880
rect 10419 41020 10561 41021
rect 10419 40860 10420 41020
rect 10560 40860 10561 41020
rect 13359 40940 13360 41040
rect 13520 40940 13521 41040
rect 16280 41021 16460 43819
rect 18830 42661 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 22199 44520 22321 44521
rect 22199 44400 22200 44520
rect 22320 44400 22321 44520
rect 22199 44399 22321 44400
rect 19240 44281 19400 44300
rect 19240 44280 19401 44281
rect 19240 44120 19260 44280
rect 19400 44120 19401 44280
rect 19240 44119 19401 44120
rect 18799 42660 18901 42661
rect 18799 42540 18800 42660
rect 18900 42540 18901 42660
rect 18799 42539 18901 42540
rect 18830 42530 18890 42539
rect 19240 41041 19400 44119
rect 13359 40939 13521 40940
rect 16279 41020 16460 41021
rect 10419 40859 10561 40860
rect 16279 40840 16280 41020
rect 16440 40840 16460 41020
rect 19239 41040 19401 41041
rect 19239 40900 19240 41040
rect 19400 40900 19401 41040
rect 22200 41021 22320 44399
rect 23798 43081 23858 45152
rect 24350 43341 24410 45152
rect 24902 43641 24962 45152
rect 25140 44761 25260 44780
rect 25139 44760 25261 44761
rect 25139 44660 25140 44760
rect 25260 44660 25261 44760
rect 25139 44659 25261 44660
rect 24839 43640 24981 43641
rect 24839 43500 24840 43640
rect 24980 43500 24981 43640
rect 24839 43499 24981 43500
rect 24902 43490 24962 43499
rect 24319 43340 24441 43341
rect 24319 43200 24320 43340
rect 24440 43200 24441 43340
rect 24319 43199 24441 43200
rect 24350 43170 24410 43199
rect 23739 43080 23901 43081
rect 23739 42920 23740 43080
rect 23900 42920 23901 43080
rect 23739 42919 23901 42920
rect 23798 42910 23858 42919
rect 22199 41020 22321 41021
rect 22199 40920 22200 41020
rect 22320 40920 22321 41020
rect 25140 40981 25260 44659
rect 25454 43981 25514 45152
rect 26006 44261 26066 45152
rect 26558 44521 26618 45152
rect 27110 44761 27170 45152
rect 27662 44761 27722 45152
rect 28214 44890 28274 45152
rect 28214 44830 28540 44890
rect 27079 44760 27181 44761
rect 27079 44640 27080 44760
rect 27180 44640 27181 44760
rect 27079 44639 27181 44640
rect 27619 44760 27761 44761
rect 27619 44640 27620 44760
rect 27760 44640 27761 44760
rect 27619 44639 27761 44640
rect 28099 44760 28201 44761
rect 28099 44640 28100 44760
rect 28200 44640 28201 44760
rect 28099 44639 28201 44640
rect 26539 44520 26621 44521
rect 26539 44420 26540 44520
rect 26620 44420 26621 44520
rect 26539 44419 26621 44420
rect 26558 44410 26618 44419
rect 25979 44260 26081 44261
rect 25979 44140 25980 44260
rect 26080 44140 26081 44260
rect 25979 44139 26081 44140
rect 26006 44130 26066 44139
rect 25419 43980 25541 43981
rect 25419 43820 25420 43980
rect 25540 43820 25541 43980
rect 25419 43819 25541 43820
rect 25454 43810 25514 43819
rect 28120 41021 28197 44639
rect 28420 42261 28540 44830
rect 28419 42260 28541 42261
rect 28419 42140 28420 42260
rect 28540 42140 28541 42260
rect 28419 42139 28541 42140
rect 28766 41921 28826 45152
rect 29318 44952 29378 45152
rect 28719 41920 28861 41921
rect 28719 41760 28720 41920
rect 28860 41760 28861 41920
rect 28719 41759 28861 41760
rect 29520 41900 29720 41920
rect 28766 41750 28826 41759
rect 29520 41720 29540 41900
rect 29700 41720 29720 41900
rect 28079 41020 28221 41021
rect 22199 40919 22321 40920
rect 25139 40980 25261 40981
rect 19239 40899 19401 40900
rect 25139 40880 25140 40980
rect 25260 40880 25261 40980
rect 28079 40920 28080 41020
rect 28220 40920 28221 41020
rect 28079 40919 28221 40920
rect 25139 40879 25261 40880
rect 25140 40840 25260 40879
rect 16279 40839 16460 40840
rect 16280 40820 16460 40839
rect 5839 36740 6001 36741
rect 5839 36600 5840 36740
rect 6000 36600 6001 36740
rect 5839 36599 6001 36600
rect 5840 36580 6000 36599
rect 5459 28860 5621 28861
rect 5459 28720 5460 28860
rect 5620 28720 5621 28860
rect 5459 28719 5621 28720
rect 5460 28700 5620 28719
rect 5059 20960 5221 20961
rect 5059 20840 5060 20960
rect 5220 20840 5221 20960
rect 5059 20839 5221 20840
rect 5061 20821 5220 20839
rect 25280 17421 25460 17740
rect 25279 17420 25461 17421
rect 25279 17280 25280 17420
rect 25460 17280 25461 17420
rect 25279 17279 25461 17280
rect 25980 17160 26140 17680
rect 25980 17000 26000 17160
rect 26120 17000 26140 17160
rect 25999 16999 26121 17000
rect 4599 16640 4750 16641
rect 4599 16500 4600 16640
rect 4720 16500 4750 16640
rect 4599 16499 4750 16500
rect 4610 16490 4750 16499
rect 15730 16620 15870 16630
rect 15730 16480 15740 16620
rect 15860 16480 15870 16620
rect 15730 7740 15870 16480
rect 29520 16260 29720 41720
rect 29520 16080 29540 16260
rect 29700 16080 29720 16260
rect 29520 16060 29720 16080
rect 15730 7600 15740 7740
rect 15860 7600 15870 7740
rect 15730 7550 15870 7600
rect 800 5940 880 6180
rect 1160 5940 1200 6180
rect 800 5320 1200 5940
rect 800 5100 920 5320
rect 1140 5100 1200 5320
rect 800 4900 1200 5100
rect 800 4620 840 4900
rect 1140 4620 1200 4900
rect 800 1000 1200 4620
rect 30362 4141 30542 4150
rect 30339 4140 30542 4141
rect 30339 3960 30340 4140
rect 30520 3960 30542 4140
rect 30339 3959 30542 3960
rect 26499 3840 26681 3841
rect 26499 3830 26500 3840
rect 26498 3660 26500 3830
rect 26680 3660 26681 3840
rect 26498 3659 26681 3660
rect 22634 3181 22814 3190
rect 22619 3180 22821 3181
rect 22619 3000 22620 3180
rect 22820 3000 22821 3180
rect 22619 2999 22821 3000
rect 18770 2701 18950 2710
rect 18759 2700 18950 2701
rect 18759 2540 18760 2700
rect 18940 2540 18950 2700
rect 18759 2539 18950 2540
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 2539
rect 22634 0 22814 2999
rect 26498 0 26678 3659
rect 30362 0 30542 3959
<< comment >>
rect 5840 17240 5860 17260
use buffer  buffer_0 /foss/designs/tt10-temp-sensor-clock-divider/mag/temp-sensor/buffer/mag
timestamp 1707919911
transform 1 0 6460 0 1 7280
box 900 -1720 7760 5820
use clock_divider  clock_divider_0
timestamp 1738624466
transform -1 0 29860 0 1 17024
box 514 496 24000 24000
use sensor  sensor_0 /foss/designs/tt10-temp-sensor-clock-divider/mag/temp-sensor/sensor/mag
timestamp 1699935153
transform 1 0 2960 0 1 8940
box -660 -2500 3580 3000
use sigma-delta  sigma-delta_0 /foss/designs/tt10-temp-sensor-clock-divider/mag/temp-sensor/sigma-delta_modulator/mag
timestamp 1729283034
transform 1 0 19080 0 1 6520
box -3180 -520 12140 5420
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
