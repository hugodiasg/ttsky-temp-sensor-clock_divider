magic
tech sky130A
magscale 1 2
timestamp 1700703435
<< metal4 >>
rect -2349 3039 2349 3080
rect -2349 -3039 2093 3039
rect 2329 -3039 2349 3039
rect -2349 -3080 2349 -3039
<< via4 >>
rect 2093 -3039 2329 3039
<< mimcap2 >>
rect -2269 2960 1731 3000
rect -2269 -2960 -2229 2960
rect 1691 -2960 1731 2960
rect -2269 -3000 1731 -2960
<< mimcap2contact >>
rect -2229 -2960 1691 2960
<< metal5 >>
rect 2051 3039 2371 3081
rect -2253 2960 1715 2984
rect -2253 -2960 -2229 2960
rect 1691 -2960 1715 2960
rect -2253 -2984 1715 -2960
rect 2051 -3039 2093 3039
rect 2329 -3039 2371 3039
rect 2051 -3081 2371 -3039
<< properties >>
string FIXED_BBOX -2349 -3080 1811 3080
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 20 l 30 val 1.219k carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
