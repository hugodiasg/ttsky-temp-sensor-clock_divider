magic
tech sky130A
magscale 1 2
timestamp 1700747285
<< nmos >>
rect -12087 -150 -6087 150
rect -6029 -150 -29 150
rect 29 -150 6029 150
rect 6087 -150 12087 150
<< ndiff >>
rect -12145 138 -12087 150
rect -12145 -138 -12133 138
rect -12099 -138 -12087 138
rect -12145 -150 -12087 -138
rect -6087 138 -6029 150
rect -6087 -138 -6075 138
rect -6041 -138 -6029 138
rect -6087 -150 -6029 -138
rect -29 138 29 150
rect -29 -138 -17 138
rect 17 -138 29 138
rect -29 -150 29 -138
rect 6029 138 6087 150
rect 6029 -138 6041 138
rect 6075 -138 6087 138
rect 6029 -150 6087 -138
rect 12087 138 12145 150
rect 12087 -138 12099 138
rect 12133 -138 12145 138
rect 12087 -150 12145 -138
<< ndiffc >>
rect -12133 -138 -12099 138
rect -6075 -138 -6041 138
rect -17 -138 17 138
rect 6041 -138 6075 138
rect 12099 -138 12133 138
<< poly >>
rect -12087 222 -6087 238
rect -12087 188 -12071 222
rect -6103 188 -6087 222
rect -12087 150 -6087 188
rect -6029 222 -29 238
rect -6029 188 -6013 222
rect -45 188 -29 222
rect -6029 150 -29 188
rect 29 222 6029 238
rect 29 188 45 222
rect 6013 188 6029 222
rect 29 150 6029 188
rect 6087 222 12087 238
rect 6087 188 6103 222
rect 12071 188 12087 222
rect 6087 150 12087 188
rect -12087 -188 -6087 -150
rect -12087 -222 -12071 -188
rect -6103 -222 -6087 -188
rect -12087 -238 -6087 -222
rect -6029 -188 -29 -150
rect -6029 -222 -6013 -188
rect -45 -222 -29 -188
rect -6029 -238 -29 -222
rect 29 -188 6029 -150
rect 29 -222 45 -188
rect 6013 -222 6029 -188
rect 29 -238 6029 -222
rect 6087 -188 12087 -150
rect 6087 -222 6103 -188
rect 12071 -222 12087 -188
rect 6087 -238 12087 -222
<< polycont >>
rect -12071 188 -6103 222
rect -6013 188 -45 222
rect 45 188 6013 222
rect 6103 188 12071 222
rect -12071 -222 -6103 -188
rect -6013 -222 -45 -188
rect 45 -222 6013 -188
rect 6103 -222 12071 -188
<< locali >>
rect -12087 188 -12071 222
rect -6103 188 -6087 222
rect -6029 188 -6013 222
rect -45 188 -29 222
rect 29 188 45 222
rect 6013 188 6029 222
rect 6087 188 6103 222
rect 12071 188 12087 222
rect -12133 138 -12099 154
rect -12133 -154 -12099 -138
rect -6075 138 -6041 154
rect -6075 -154 -6041 -138
rect -17 138 17 154
rect -17 -154 17 -138
rect 6041 138 6075 154
rect 6041 -154 6075 -138
rect 12099 138 12133 154
rect 12099 -154 12133 -138
rect -12087 -222 -12071 -188
rect -6103 -222 -6087 -188
rect -6029 -222 -6013 -188
rect -45 -222 -29 -188
rect 29 -222 45 -188
rect 6013 -222 6029 -188
rect 6087 -222 6103 -188
rect 12071 -222 12087 -188
<< viali >>
rect -12071 188 -6103 222
rect -6013 188 -45 222
rect 45 188 6013 222
rect 6103 188 12071 222
rect -12133 -121 -12099 17
rect -6075 -17 -6041 121
rect -17 -121 17 17
rect 6041 -17 6075 121
rect 12099 -121 12133 17
rect -12071 -222 -6103 -188
rect -6013 -222 -45 -188
rect 45 -222 6013 -188
rect 6103 -222 12071 -188
<< metal1 >>
rect -12083 222 -6091 228
rect -12083 188 -12071 222
rect -6103 188 -6091 222
rect -12083 182 -6091 188
rect -6025 222 -33 228
rect -6025 188 -6013 222
rect -45 188 -33 222
rect -6025 182 -33 188
rect 33 222 6025 228
rect 33 188 45 222
rect 6013 188 6025 222
rect 33 182 6025 188
rect 6091 222 12083 228
rect 6091 188 6103 222
rect 12071 188 12083 222
rect 6091 182 12083 188
rect -6081 121 -6035 133
rect -12139 17 -12093 29
rect -12139 -121 -12133 17
rect -12099 -121 -12093 17
rect -6081 -17 -6075 121
rect -6041 -17 -6035 121
rect 6035 121 6081 133
rect -6081 -29 -6035 -17
rect -23 17 23 29
rect -12139 -133 -12093 -121
rect -23 -121 -17 17
rect 17 -121 23 17
rect 6035 -17 6041 121
rect 6075 -17 6081 121
rect 6035 -29 6081 -17
rect 12093 17 12139 29
rect -23 -133 23 -121
rect 12093 -121 12099 17
rect 12133 -121 12139 17
rect 12093 -133 12139 -121
rect -12083 -188 -6091 -182
rect -12083 -222 -12071 -188
rect -6103 -222 -6091 -188
rect -12083 -228 -6091 -222
rect -6025 -188 -33 -182
rect -6025 -222 -6013 -188
rect -45 -222 -33 -188
rect -6025 -228 -33 -222
rect 33 -188 6025 -182
rect 33 -222 45 -188
rect 6013 -222 6025 -188
rect 33 -228 6025 -222
rect 6091 -188 12083 -182
rect 6091 -222 6103 -188
rect 12071 -222 12083 -188
rect 6091 -228 12083 -222
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.5 l 30 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc -50 viadrn +50 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
